////////////////////////////////////////////////////////////////////////////////
//(c) Copyright 2013 Mobiveil, Inc. All rights reserved
//
// File    :  srio_ll_atomic_dec_test.sv
// Project :  srio vip
// Purpose : Atomic  decrement test 
// Author  :  Mobiveil
//
// Test for Atomic  decrement.
//
////////////////////////////////////////////////////////////////////////////////

class srio_ll_atomic_dec_test extends srio_base_test;

  `uvm_component_utils(srio_ll_atomic_dec_test)

  srio_ll_atomic_dec_seq atomic_dec_seq;

    
  function new(string name, uvm_component parent=null);
    super.new(name, parent);
  endfunction

    task run_phase( uvm_phase phase );
    super.run_phase(phase);
    atomic_dec_seq = srio_ll_atomic_dec_seq::type_id::create("atomic_dec_seq");

      phase.raise_objection( this );
     atomic_dec_seq.start( env1.e_virtual_sequencer);
     
  #20000ns;
    phase.drop_objection(this);
    
  endtask

  
endclass


