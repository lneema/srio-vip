////////////////////////////////////////////////////////////////////////////////
//(c) Copyright 2013 Mobiveil, Inc. All rights reserved
//
// File    :  srio_tl_variables.sv
// Project :  srio vip
// Purpose :  Transport Layer Variables
// Author  :  Mobiveil
//
// TL Variables
//
//////////////////////////////////////////////////////////////////////////////// 
typedef class srio_tl_sequencer;                                                            
typedef class srio_tl_bfm;                                                                  
typedef class srio_tl_config;                                                               
typedef class srio_tl_generator;                                                              
typedef class srio_tl_receiver;                                                               
typedef class srio_tl_monitor;
typedef class srio_tl_txrx_monitor;
