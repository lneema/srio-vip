
////////////////////////////////////////////////////////////////////////////////
//(c) Copyright 2013 Mobiveil, Inc. All rights reserved
//
// File    : srio_pl_random_acc_gen_kind_test .sv
// Project :  srio vip
// Purpose :  NREAD
// Author  :  Mobiveil
//
// 1. Set PL_RANDOM acc gen kind value..now the ackid value generate in random delay.
// 2.Test for NREAD request class
//
////////////////////////////////////////////////////////////////////////////////

class srio_pl_random_acc_gen_kind_test extends srio_base_test;

  `uvm_component_utils(srio_pl_random_acc_gen_kind_test)

  srio_ll_nread_req_seq nread_req_seq;

    
  function new(string name, uvm_component parent=null);
    super.new(name, parent);
  endfunction

    task run_phase( uvm_phase phase );
    super.run_phase(phase);
    env_config2.pl_config.pkt_acc_gen_kind = PL_RANDOM; 
    nread_req_seq = srio_ll_nread_req_seq::type_id::create("nread_req_seq");

     phase.raise_objection( this );
      nread_req_seq.start( env1.e_virtual_sequencer);
      #2000ns;
 
    phase.drop_objection(this);
    
  endtask

  
endclass


