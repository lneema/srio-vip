////////////////////////////////////////////////////////////////////////////////////////////////
//(c) Copyright 2013 Mobiveil, Inc. All rights reserved
//
// File       :  srio_pl_lane_handler.sv
// Project    :  srio vip
// Purpose    :  Lane handler class. It performs the following functions,
// 		 1. SIPO
// 		 2. 10b to 8b decoding / 67b to 64b decoding
// 		 3. Descramling.
// 		 4. Lane specific state machines
//		 5. IDLE2 AET, GEN3 CW training, GEN3 DME training.
// Author     :  Mobiveil
//
// Physical layer lane handler class.
//
//
//////////////////////////////////////////////////////////////////////////////////////////////////

class srio_pl_lane_handler extends uvm_component;

  /// @cond
  `uvm_component_utils(srio_pl_lane_handler)
  /// @endcond

  
  virtual srio_interface srio_if;			///< Virtual interface

  srio_env_config lh_env_config;			///< ENV Config instance

  srio_pl_config lh_config;				///< PL Config instance

  srio_pl_common_component_trans lh_trans;		///< PL monitor common transaction instance

  srio_pl_tx_rx_mon_common_trans lh_common_mon_trans;	///< Common monitor transction instance

  srio_reg_block lh_reg_model;				///< Register model instance

  // Properties
  int lane_num;						///< lane number
  int invalid_cg_cnt;					///< Invalid codegroup count after s2p_lock is set.

  srio_pl_lane_data lane_data_ins;			///< lane data instance. It contains all the information related
  srio_pl_lane_data temp_lane_data_ins;			///< lane data instance. It contains all the information related
							///< to the 10 bit serial data, its 8bit decoded value etc.

  bit rx_clk;						///< rx_clk generated from lane specific rx_clk in interface
  bit tx_clk;						///< tx_clk generated from lane specific tx_clk in interface
  bit rx_data;						///< rx data generated from lane specific rx_data in interface
  bit divide_clk;					///< divide_clk generated by locking comma character
  bit s2p_lock;						///< indicates 10-bit or 67-bit lock is acheived.

  bit [0:9] rx_pdata;					///< rx data generated from lane specific rx_data in interface
 
  bit bfm_or_mon;					///< 1 : bfm instance ; 0 : monitor instance
  bit mon_type;						///< 1 : tx_monitor ; 0 : rx_monitor
  bit report_error;					///< 1 : error ; 0 : warning

  bit dut_tx_scr_dis;					///< dut tx scrambling disable.
  bit dut_rcvr_trn_spt;					///< dut receiver trained support.
  bit dut_rcvr_trn_en;					///< dut receiver trained enable.
  bit descr_in_sync;					///< GEN2.x descrambler is in sync.
  bit [16:0] descr_lfsr;				///< lfsr used for GEN2.x descrambling.
  bit start_descr_sync;					///< Indicates GEN2.x descrambler sync can be started.
  bit descr_sync_check;					///< Indicates GEN2.x descrambler sync check is being performed.

  int M_cnt;						///< 'M' character count used for descrambler sync check.
  int cs_field_byte_cnt;				///< No. of bytes received in CS field.
  int D_after_M_cnt;					///< No. of data characters received after an 'M', to detect MDDDD.
  int descr_sync_check_cnt;				///< Descrambler sync check counter.

  bit prev_idle2_cs;					///< Previous value of idle2_cs.
  int K_counter;					///< 'K' character counter used in Sync state machine.
  int V_counter;					///< Valid character counter used in Sync state machine.
  int I_counter;					///< Invalid character counter used in Sync state machine.
  int IV_counter;					///< Invalid counter used in gen3 codeword lock state machine.
  int CW_counter;					///< Codeword counter used in gen3 codeword lock state machine.

  bit ls0_rcvr_pol_field_updated;			///< Receiver polarity. Used to update the corresponding register.

  bit check_cmd_deassertion;				///< IDLE2 AET command deassertion check enabled.
  bit check_cmd_reassertion;				///< IDLE2 AET command reassertion check enabled.
  bit cmd_reassertion_timer_done;			///< IDLE2 AET command reassertion timer completed.
  bit idle2_cs_field_started;				///< Indicates IDLE2 cs field is being received.
  int idle2_aet_cmd_cnt;				///< IDLE2 AET command count to check multiple command assertion in a single CS field.
  int idle2_cs_fld_method_char_cnt;			///< Characters count to collect complete CS field.

  bit idle2_value_changed;				///< Bit used to update IDLE2 related register field.
  bit [0:2] idle2_cs_marker_port_width;			///< Variable used to update IDLE2 related register field.
  bit [0:3] idle2_cs_marker_lane_number;		///< Variable used to update IDLE2 related register field.

  bit [0:31] lane_status_1_reg_val;			///< Variable used to update IDLE2 related register field.

  srio_pl_rcvd_cs_field_data lane_cs_fld_data_ins;	///< Instances of srio_pl_rcvd_cs_field_data. Used in IDLE2 AET checks.
  srio_pl_rcvd_cs_field_data prev_lane_cs_fld_data_ins;
  srio_pl_rcvd_cs_field_data bkp_lane_cs_fld_data_ins;

  sync_sm_states prev_sync_state, current_sync_state;	///< Indicates current and previous sync states.
  sync_sm_states current_sync_state_q[$];		///< current sync state queue for FC to hit intermediate states.

  // GEN3.0 variables

  bit [0:66] gen3_rx_pdata;				///< GEN3.0 rx parallel data generated from lane specific rx_data in interface
  bit [0:66] gen3_rx_pdata_tmp;				///< GEN3.0 rx parallel data generated from lane specific rx_data in interface

  bit [0:57] gen3_descr_lfsr;				///< GEN3.0 descrambler LFSR.
  bit [0:57] temp_gen3_descr_lfsr;			///< Temporary variable for GEN3.0 descrambler LFSR.

  bit [57:0] reversed_gen3_descr_lfsr;			///< Reversed version of GEN3.0 descrambler LFSR.
  bit [57:0] reversed_temp_gen3_descr_lfsr;		///< Reversed version of GEN3.0 temp descrambler LFSR.

  bit [0:57] gen3_shifted_lfsr;				///< Holds the shifted value of GEN3.0 Descrambler LFSR

  int descr_seed_cntl_cw_cnt;				///< Used to detect the occurance of descr-seed control cw in the descr-seed ordered sequence.
  int sync1_state_ui_cnt;				///< Unit interval count used in GEN3.0 sync state machine.

  bit [0:63] prev_status_cntl_cw;			///< Holds the first status control control codeword of status/control ordered sequence.

  bit sync_sm_descr_sync;				///< Indicates descrambler is in sync. Used in GEN3.0 sync state machine.
  bit sync_sm_descr_err;				///< Indicates descrambler error. Used in GEN3.0 sync state machine.

  int lh_status_cntl_cw_cnt;				///< Used to detect the occurance of stat-cntl control cw in the stat-cntl ordered sequence.
  int lh_descr_seed_cw_cnt;				///< Used to detect the occurance of descr-seed control cw in the descr-seed ordered sequence.
  int lh_skip_os_cw_cnt;				///< Used to detect control CWs in the SKIP ordered sequence.

  bit trigger_os_check_methods;				///< Indicates checking of ordered sequence can be started.

  bit gen3_cmd_deassertion_timer_done;			///< Indicates GEN3.0 training command deassertion timer is completed.

  bit dme_frame_divide_clk;				///< divide_clk generated by locking DME frame marker
  bit dme_frame_s2p_lock;				///< indicates 67-bit lock is acheived for DME frame.

  bit [0:4383] complete_dme_frame;			///< Holds a complete DME frame at a time.

  int frame_bit_count;					///< Counts the number of DME frame bits received.
  int temp_frame_bit_count;				///< Temp variable used for frame_bit_count.
  int remaining_bits_in_prev_frame;			///< Indicates the remaining bits in previous frame.
  int temp_remaining_bits;				///< Temp variable used for remaining_bits_in_prev_frame.

  bit frame_offset;					///< Indicates a complete frame is received.
  bit frame_offset_achieved;				///< Temp variable used for frame_offset as it'll be cleared in the frame-lock state machine.
  bit gen3_parallel_mode_frame_received;		///< Indicates frame is locked in parallel mode.
  bit parallel_slide_mode=0;

  bit new_marker;					///< Indicates new frame marker is received.

  bit [0:31] frame_marker_data;				///< Contains the value of frame marker received.
  
  int good_markers;					///< Indicates the count of good frame markers received.
  int bad_markers;					///< Indicates the count of bad frame markers received.

  bit slip_done;					///< Indicates that dme_frame_s2p_lock is cleared after set, 
							///< and serial data is shifted to next position to check the frame position.

  bit [0:255] dme_coeff_update_status_field;		///< Holds a complete control channel of a DME frame.
  bit [0:31] decoded_dme_data;				///< Holds the decoded control channel of a DME frame.
  bit [15:0] decoded_dme_coeff_update_field;		///< Contains the decoded coefficient update field of a DME frame.
  bit [15:0] decoded_dme_status_field;			///< Contains the decoded status field of a DME frame.

  int c0_preset_value;					///< Preset value of c0 tap used in long-run training.
  int c0_init_value;					///< Initialize value of c0 tap used in long-run training.
  int c0_max_limit;					///< Maximum limit for c0 tap coefficient value used in long-run training.
  int c0_min_limit;					///< Minimum limit for c0 tap coefficient value used in long-run training.

  int cp1_preset_value;					///< Preset value of cp1 tap used in long-run training.
  int cp1_init_value;    				///< Initialize value of cp1 tap used in long-run training.
  int cp1_max_limit;     				///< Maximum limit for cp1 tap coefficient value used in long-run training.
  int cp1_min_limit;     				///< Minimum limit for cp1 tap coefficient value used in long-run training.

  int cn1_preset_value;					///< Preset value of cn1 tap used in long-run training.
  int cn1_init_value;    				///< Initialize value of cn1 tap used in long-run training.
  int cn1_max_limit;     				///< Maximum limit for cn1 tap coefficient value used in long-run training.
  int cn1_min_limit;     				///< Minimum limit for cn1 tap coefficient value used in long-run training.

  int new_c0_coeff;					///< New c0 tap coefficient value.
  int new_cp1_coeff;					///< New cp1 tap coefficient value.
  int new_cn1_coeff;					///< New cn1 tap coefficient value.

  bit [0:31] ls2_reg_val;				///< Holds the Lane N status 2 register update value.
  bit [0:31] ls3_reg_val;				///< Holds the Lane N status 3 register update value.

  bit [0:22] bip23_value;				///< Holds the expected BIP23 value.
  bit [0:22] temp_bip23_value;				///< Holds the BIP23 value calculated from the current codeword.
  bit lc_after_cw_lock_detected;			///< Indicates first lane check control codeword is detected after codeword lock.
  int note_bit_1=67;                                    ///< Marker to hold the slip information on parallel data
  int note_bit_2=66;                                    ///< Marker to hold the slip information on parallel data
  int note_bit_3=67;                                    ///< Marker to hold the slip information on parallel data
  bit [0:66] sixty_seven_bit_data;
  bit [0:66] sixty_seven_bit_data_reg;
  bit [0:66] sixty_seven_bit_data_tmp=0;
  cw_lock_sm_states prev_cw_lock_state, current_cw_lock_state;		///< Indicates current and previous CW lock state.
  cw_lock_sm_states current_cw_lock_state_q[$];				///< current CW lock state queue for FC to hit intermediate states.

  srio_pl_gen3_lane_train_data gen3_train_data_ins;			///< srio_pl_gen3_lane_train_data instances used for long-run training checks.
  srio_pl_gen3_lane_train_data bkp_gen3_train_data_ins;

  link_train_sm_states prev_cw_train_state, current_cw_train_state;	///< current and previous short-run training states.
  link_train_sm_states prev_dme_train_state, current_dme_train_state;	///< current and previous long-run training states.
  link_train_sm_states current_cw_train_state_q[$];                     ///< current and previous short-run training states queue ti hit FC
  link_train_sm_states current_dme_train_state_q[$];                    ///< current and previous long-run training states queue ti hit FC

  frame_lock_sm_states prev_frame_lock_state, current_frame_lock_state;	///< current and previous frame lock states.

  dme_training_coeff_update_states prev_c0_coeff_update_state, current_c0_coeff_update_state;	///< current and previous c0 tap coefficient update states.
  dme_training_coeff_update_states prev_cp1_coeff_update_state, current_cp1_coeff_update_state;	///< current and previous cp1 tap coefficient update states.
  dme_training_coeff_update_states prev_cn1_coeff_update_state, current_cn1_coeff_update_state;	///< current and previous cn1 tap coefficient update states.
  frame_lock_sm_states current_frame_lock_state_q[$];
  dme_training_coeff_update_states current_c0_coeff_update_state_q[$];
  dme_training_coeff_update_states current_cp1_coeff_update_state_q[$];
  dme_training_coeff_update_states current_cn1_coeff_update_state_q[$];

  uvm_reg_field reqd_field_name[string];	///< Associative array to get respective field name from register_update_method.

  // Events
  uvm_event srio_rx_lane_event;			///< Event used to pass the lane data to higher level component.

  event start_100us_cmd_timer;			///< Triggers the 100us command timer. Used in short-run training checks.
  
  // Callback register
  `uvm_register_cb(srio_pl_lane_handler, srio_pl_callback)	///< Registering PL callback

  // Methods
  extern function new(string name = "srio_pl_lane_handler", uvm_component parent = null);
  extern task run_phase(uvm_phase phase);
  
  extern virtual task rx_clk_data_gen();
  extern virtual task ser2par();
  extern virtual task tenb_8b_decode();
  extern virtual task calc_curr_rd(input int data);
  extern virtual task init_lfsr();
  extern virtual task shift_descr_lfsr();
  extern virtual task data_descramble();
  extern virtual task lane_sync_sm();
  extern virtual task lane_ready_gen();
  extern virtual task collect_idle2_csfield();
  extern virtual task idle2_aet_method();
  extern virtual task idle2_aet_checks();
  extern virtual task idle2_aet_timer_method();
  extern virtual task set_receiver_trained();
  extern virtual task comma_char_freq_check();

  extern virtual task update_ls0_lane_num_field();
  extern virtual task update_ls0_8b_10b_dec_err_field();
  extern virtual task update_ls0_rcvr_pol_field();
  extern virtual task update_other_ls0_fields();
  extern virtual task update_ls1_reg();

  // GEN3.0 methods

  extern virtual task sixty_sevenb_sixty_fourb_decode();
  extern virtual task gen3_data_descramble();
  extern virtual task status_cntl_os_check_method();
  extern virtual task descr_seed_os_check_method();
  extern virtual task skip_os_check_method();
  extern virtual task skip_marker_cw_fixed_value_check();
  extern virtual task skip_cw_fixed_value_check();
  extern virtual task gen3_cw_training_method();
  extern virtual task gen3_training_checks();
  extern virtual task gen3_cw_training_cmd_timer_method();
  extern virtual task shift_gen3_descr_lfsr(int shift_count, bit [0:57] gen3_lfsr); // task with ref argument needs to be automatic
  extern virtual task cw_lock_sm();
  extern virtual task gen3_lane_sync_sm();
  extern virtual task gen3_cw_training_sm();
  extern virtual task gen3_train_timer();
  extern virtual task gen3_keep_alive_timer_method();

  extern virtual task gen3_frame_lock_sm();
  extern virtual task gen3_dme_training_sm();
  extern virtual task gen3_dme_training_commands_decode();
  extern virtual task gen3_dme_decode(bit [0:255] dme_data);
  extern virtual task dme_wait_timer_method();

  extern virtual task gen3_c0_coeff_update_sm();
  extern virtual task gen3_cp1_coeff_update_sm();
  extern virtual task gen3_cn1_coeff_update_sm();
  extern virtual task lc_cw_bip_calc_method();

  extern virtual task update_ls1_idle3_training_type(bit [2:0] training_type_val);
  extern virtual task update_ls1_idle3_dme_training_state();
  extern virtual task update_ls1_idle3_cw_training_state();
  extern virtual task update_ls1_idle3_cw_retraining_state();
  extern virtual task update_ls2_reg();
  extern virtual task update_ls3_reg();

  extern virtual task update_error_detect_csr(string csr_field_name);

  extern virtual task automatic register_update_method(string reg_name, string field_name, int offset, string reg_ins, output uvm_reg_field out_field_name);

  // Callback related methods

  virtual task srio_pl_cg_received_lane0(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane1(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane2(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane3(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane4(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane5(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane6(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane7(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane8(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane9(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane10(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane11(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane12(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane13(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane14(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_cg_received_lane15(ref srio_pl_lane_data rx_srio_cg, srio_env_config lh_env_config);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane0(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane1(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane2(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane3(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane4(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane5(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane6(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane7(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane8(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane9(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane10(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane11(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane12(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane13(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane14(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 
  
  virtual task srio_pl_aet_cs_received_lane15(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
  endtask 

  /*task temp_8b_data_to_if();

    forever begin //{

      if (lane_num == 0)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_0 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 1)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_1 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 2)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_2 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 3)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_3 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 4)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_4 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 5)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_5 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 6)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_6 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 7)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_7 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 8)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_8 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 9)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_9 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 10)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_10 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 11)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_11 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 12)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_12 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 13)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_13 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 14)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_14 = lane_data_ins.brc3_cw;
      end //}
      else if (lane_num == 15)
      begin //{
        @(lane_data_ins.brc3_cw)
          srio_if.env_rxdata_15 = lane_data_ins.brc3_cw;
      end //}

    end //}

  endtask

  task temp_8b_cntl_to_if();

    forever begin //{

      if (lane_num == 0)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_0 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 1)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_1 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 2)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_2 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 3)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_3 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 4)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_4 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 5)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_5 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 6)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_6 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 7)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_7 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 8)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_8 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 9)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_9 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 10)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_10 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 11)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_11 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 12)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_12 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 13)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_13 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 14)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_14 = lane_data_ins.cntl;
      end //}
      else if (lane_num == 15)
      begin //{
        @(lane_data_ins.cntl)
          srio_if.env_rxcntl_15 = lane_data_ins.cntl;
      end //}

    end //}

  endtask*/

endclass


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : New
/// Description : Constructor method for srio_pl_lane_handler class.
///////////////////////////////////////////////////////////////////////////////////////////////
function srio_pl_lane_handler::new(string name="srio_pl_lane_handler", uvm_component parent=null);
  super.new(name, parent);
  lane_data_ins = new();
  lane_data_ins.curr_rd = NEG;
endfunction : new



///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : run_phase
/// Description : run_phase method of srio_pl_lane_handler class.
/// It triggers all the methods within the class which needs to be run forever.
/// It also registers the callback for uvm_error demote logic.
///////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::run_phase(uvm_phase phase);

  err_demoter pl_lh_err_demoter = new();
  pl_lh_err_demoter.en_err_demote = !report_error;
  uvm_report_cb::add(this, pl_lh_err_demoter);

  if (~bfm_or_mon)
  begin //{

    lh_common_mon_trans.idle2_aet_cmd_outstanding[mon_type][lane_num] = 1;
    lh_common_mon_trans.idle2_aet_cmd_outstanding[mon_type][lane_num] = 0;

    lh_common_mon_trans.idle2_aet_ack_nack_rcvd[mon_type][lane_num] = 1;
    lh_common_mon_trans.idle2_aet_ack_nack_rcvd[mon_type][lane_num] = 0;

    lh_common_mon_trans.command_deasserted[mon_type][lane_num] = 1;
    lh_common_mon_trans.command_deasserted[mon_type][lane_num] = 0;

  end //}

  fork

    rx_clk_data_gen();
    ser2par();
    lane_ready_gen();
    set_receiver_trained();

    if (~bfm_or_mon)
      comma_char_freq_check();

    if (lh_env_config.srio_mode != SRIO_GEN30)
    begin //{

      fork
        lane_sync_sm();
        collect_idle2_csfield();
        if (~bfm_or_mon)
          idle2_aet_timer_method();
        //if (bfm_or_mon)
        //  temp_8b_data_to_if();
        //if (bfm_or_mon)
        //  temp_8b_cntl_to_if();
        if (~bfm_or_mon)
          update_ls0_8b_10b_dec_err_field();
      join_none

    end //}
    else
    begin //{
      fork

        cw_lock_sm();
        gen3_lane_sync_sm();
        gen3_cw_training_sm();
        gen3_cw_training_cmd_timer_method();
        gen3_train_timer();
        gen3_keep_alive_timer_method();

	if (lh_config.brc3_training_mode)
	  gen3_frame_lock_sm();

	if (lh_config.brc3_training_mode)
	  gen3_dme_training_sm();

	if (~bfm_or_mon && lh_config.brc3_training_mode)
	  dme_wait_timer_method();

	if (lh_config.brc3_training_mode)
	  gen3_dme_training_commands_decode();

	if (lh_config.brc3_training_mode)
	  gen3_c0_coeff_update_sm();

	if (lh_config.brc3_training_mode)
	  gen3_cp1_coeff_update_sm();

	if (lh_config.brc3_training_mode)
	  gen3_cn1_coeff_update_sm();

      join_none
    end //}

  join_none

endtask : run_phase



///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : rx_clk_data_gen
/// Description : This method takes a local copy of the clock and data declared in the interface,
/// based on the srio_interface_mode, bfm_or_mon and mon_type.
///////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::rx_clk_data_gen();
 int slice=0;
 int lsb=0;
  if (lh_env_config.srio_interface_mode == SRIO_SERIAL)
  begin //{

    fork //{

        begin //{
         forever
          begin //{
             @(srio_if.tx_sclk[lane_num]);
             tx_clk = srio_if.tx_sclk[lane_num];
          end //}
        end //}
      begin //{

        forever
        begin //{

	  @(srio_if.rx_sclk[lane_num]);
	  rx_clk = srio_if.rx_sclk[lane_num];

        end //}

      end //}


      begin //{

        forever
        begin //{

          if (bfm_or_mon)
          begin //{

	    @(srio_if.rxp[lane_num]);
	    rx_data = srio_if.rxp[lane_num];

          end //}
          else if (~mon_type)  // tx_mon or rx_mon
          begin //{

	    @(srio_if.rxp[lane_num]);
	    rx_data = srio_if.rxp[lane_num];

          end //}
          else
          begin //{

	    @(srio_if.txp[lane_num]);
	    rx_data = srio_if.txp[lane_num];

          end //}

        end //}

      end //}

    join //}

  end //}
  else if (lh_env_config.srio_interface_mode == SRIO_PARALLEL)
  begin //{

    fork //{
        begin //{
         forever
          begin //{
             @(srio_if.tx_pclk[lane_num]);
             tx_clk = srio_if.tx_pclk[lane_num];

          if(mon_type)
	  divide_clk = tx_clk;

	  if (lh_env_config.srio_mode == SRIO_GEN30 && lh_config.brc3_training_mode && mon_type)
	    dme_frame_divide_clk = tx_clk;
          end //}
        end //}

      begin //{

        forever
        begin //{

	  @(srio_if.rx_pclk[lane_num]);
	  rx_clk = srio_if.rx_pclk[lane_num];

          if(~mon_type)
	  divide_clk = rx_clk;

	  if (lh_env_config.srio_mode == SRIO_GEN30 && lh_config.brc3_training_mode && ~mon_type)
	    dme_frame_divide_clk = rx_clk;

        end //}

      end //}


      begin //{

        forever
        begin //{

          if (bfm_or_mon)
          begin //{

	    if (lh_env_config.srio_mode != SRIO_GEN30)
	    begin //{
	      @(srio_if.rx_pdata[lane_num]);
	      rx_pdata = srio_if.rx_pdata[lane_num];
	    end //}
	    else
	    begin //{
	      //@(srio_if.gen3_rx_pdata[lane_num]);
         	@(posedge srio_if.rx_pclk[lane_num]);
                 begin//{
                  if(~lh_config.parallel_dme_slip_adj_en)
	           gen3_rx_pdata = srio_if.gen3_rx_pdata[lane_num];
                  else
	           begin //{
	            gen3_rx_pdata_tmp = srio_if.gen3_rx_pdata[lane_num];
                    if(~parallel_slide_mode || (note_bit_2==0))
                     begin//{
                      gen3_rx_pdata=gen3_rx_pdata_tmp;
                     end//}
                    else
                     begin//{
                      slice=67-note_bit_2;
                      lsb=0;
                      for(int i=slice;i<67;i++)
                       begin//{
                       gen3_rx_pdata[i]=gen3_rx_pdata_tmp[lsb];
                       lsb++;
                       end//}
                      gen3_rx_pdata_tmp=gen3_rx_pdata_tmp<<note_bit_2;
                     end//}
                   end//}
                 end//}
	    end //}

          end //}
          else if (~mon_type)  // tx_mon or rx_mon
          begin //{

	    if (lh_env_config.srio_mode != SRIO_GEN30)
	    begin //{
	      @(srio_if.rx_pdata[lane_num]);
	      rx_pdata = srio_if.rx_pdata[lane_num];
	    end //}
	    else
	    begin //{
	      //@(srio_if.gen3_rx_pdata[lane_num]);
	      @(posedge srio_if.rx_pclk[lane_num]);
               begin//{
                if(~lh_config.parallel_dme_slip_adj_en)
	         gen3_rx_pdata = srio_if.gen3_rx_pdata[lane_num];
               else
	        begin //{
	         gen3_rx_pdata_tmp = srio_if.gen3_rx_pdata[lane_num];
                 if(~parallel_slide_mode|| (note_bit_2==0))
                  begin//{
                   gen3_rx_pdata=gen3_rx_pdata_tmp;
                  end//}
                 else
                  begin//{
                   slice=67-note_bit_2;
                   lsb=0;
                   for(int i=slice;i<67;i++)
                    begin//{
                    gen3_rx_pdata[i]=gen3_rx_pdata_tmp[lsb];
                    lsb++;
                    end//}
                   gen3_rx_pdata_tmp=gen3_rx_pdata_tmp<<note_bit_2;
                  end//}
                end//}
               end//}
	    end //}

          end //}
          else
          begin //{

	    if (lh_env_config.srio_mode != SRIO_GEN30)
	    begin //{
	      @(srio_if.tx_pdata[lane_num]);
	      rx_pdata = srio_if.tx_pdata[lane_num];
	    end //}
	    else
	    begin //{
             @(posedge srio_if.tx_pclk[lane_num]);
	     // @(srio_if.gen3_tx_pdata[lane_num]);
              begin//{
               if(~lh_config.parallel_dme_slip_adj_en)
	        gen3_rx_pdata = srio_if.gen3_tx_pdata[lane_num];
               else
                begin//{
	         gen3_rx_pdata_tmp = srio_if.gen3_tx_pdata[lane_num];
                 if(~parallel_slide_mode|| (note_bit_2==0))
                  begin//{
                   gen3_rx_pdata=gen3_rx_pdata_tmp;
                  end//}
                 else
                  begin//{
                   slice=67-note_bit_2;
                   lsb=0;
                   for(int i=slice;i<67;i++)
                    begin//{
                    gen3_rx_pdata[i]=gen3_rx_pdata_tmp[lsb];
                    lsb++;
                    end//}
                   gen3_rx_pdata_tmp=gen3_rx_pdata_tmp<<note_bit_2;
                  end//}
                end//}
              end//}
	    end //}

          end //}

        end //}

      end //}

    join //}

  end //}

endtask : rx_clk_data_gen



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : ser2par
/// Description : For GEN1.3 and GEN2.x, this method performs the serial to parallel conversion,
/// based on the srio_interface_mode configured. Forms the 10-bit data and if that matches with 
/// the comma character based on the current running disparity, then  lock the 10-bit position. 
/// If the sync SM detects multiple invalid characters, then the lock mechanism is performed 
/// again. Data sampled by the SYNC sm will be decoded and descrambled data. divide_clk is also 
/// generated inside this method. divide_clk is always zero until s2p_lock is set. Once the 
/// s2p_lock is set, the divide_clk is toggled for every 5 count of ten_bit_cnt which inherently 
/// matches 5 rx_clk cycles.
/// Similarly for GEN3.0, it forms the 67-bit data code-words, generates divide-by-67 clock, decodes,
/// descrambles and keeps the data ready to be sampled by CW lock sm, frame lock sm and lane sync sm.
/// It also triggers the methods used to collect data required for adaptive equalization.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::ser2par();

  int ten_bit_cnt;
  bit [0:9] ten_bit_data;

  int sixty_seven_bit_cnt;
  int dme_frame_sixty_seven_bit_cnt;
  bit [0:66] dme_frame_sixty_seven_bit_data=0;
  bit [0:66] dme_frame_sixty_seven_bit_data_tmp=0;

  bit [0:66] brc3_frame_data;
  int slice=0;
  int lsb=0;

  forever
  begin //{

//    @(posedge rx_clk)
        if (bfm_or_mon === 0 && mon_type === 1)
           @(negedge tx_clk);
        else
          @(posedge rx_clk);
    begin //{

      if ((~s2p_lock && lh_env_config.srio_interface_mode == SRIO_SERIAL) || (~s2p_lock && lh_env_config.srio_interface_mode == SRIO_PARALLEL))
      begin //{
  //      if(~s2p_lock && lh_env_config.srio_interface_mode == SRIO_SERIAL)
	 divide_clk = 0;
	lh_trans.signal_detect[lane_num] = 0;
        note_bit_1=67;
      end //}

      if (~dme_frame_s2p_lock && lh_env_config.srio_interface_mode == SRIO_SERIAL)
      begin //{
	dme_frame_divide_clk = 0;
      end //}

      if (lh_env_config.srio_mode !== SRIO_GEN30)
      begin //{

        if (lh_env_config.srio_interface_mode == SRIO_SERIAL)
        begin //{

          ten_bit_data = ten_bit_data<<1;
          ten_bit_data[9] = rx_data;
          ten_bit_cnt++;

        end //}
        else if (lh_env_config.srio_interface_mode == SRIO_PARALLEL)
        begin //{

          ten_bit_data = rx_pdata;

        end //}

        if (lh_env_config.srio_interface_mode == SRIO_SERIAL)
        begin //{

          if (ten_bit_cnt == 10 && ~s2p_lock)
          begin //{

            if (lh_env_config.srio_mode == SRIO_GEN13)
            begin //{

              if (lane_data_ins.curr_rd == POS && ten_bit_data == 10'h305)
                s2p_lock = 1;
              else if (lane_data_ins.curr_rd == NEG && ten_bit_data == 10'hFA)
                s2p_lock = 1;
              else
                ten_bit_cnt--;

            end //}
            else if (lh_env_config.srio_mode == SRIO_GEN21 || lh_env_config.srio_mode == SRIO_GEN22)
            begin //{

              if (lane_data_ins.curr_rd == POS && (ten_bit_data == 10'h305 || ten_bit_data == 10'h306))
                s2p_lock = 1;
              else if (lane_data_ins.curr_rd == NEG && (ten_bit_data == 10'hFA || ten_bit_data == 10'hF9))
                s2p_lock = 1;
              else
                ten_bit_cnt--;

            end //}

//          `uvm_info("SRIO_LANE_HANDLER :", $sformatf("LANE NUM : %0d CHAR %0h received, CURRENT RUNNING DISPARITY is %0s", lane_num, ten_bit_data, lane_data_ins.curr_rd.name()), UVM_LOW)


          end //}

          if (ten_bit_cnt == 5 && s2p_lock)
            divide_clk = ~divide_clk;

        end //}

        if ((ten_bit_cnt == 10 && s2p_lock) || lh_env_config.srio_interface_mode == SRIO_PARALLEL)
        begin //{

//        `uvm_info("SRIO_LANE_HANDLER :", $sformatf("LANE NUM : %0d AFter s2p_lock set. CHAR %0h received, CURRENT RUNNING DISPARITY is %0s", lane_num, ten_bit_data, lane_data_ins.curr_rd.name()), UVM_LOW)

          lh_trans.signal_detect[lane_num] = 1;

          if (lh_env_config.srio_interface_mode == SRIO_SERIAL)
            ten_bit_cnt = 0;

          if (lh_trans.lane_polarity_inverted)
          begin //{
            ten_bit_data = ~ten_bit_data;
            if (~ls0_rcvr_pol_field_updated && ~bfm_or_mon)
              update_ls0_rcvr_pol_field();
          end //}

          lane_data_ins.cg = ten_bit_data;

          if (bfm_or_mon)
          begin //{

            if (lane_num == 0)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane0(lane_data_ins, lh_env_config))
            else if (lane_num == 1)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane1(lane_data_ins, lh_env_config))
            else if (lane_num == 2)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane2(lane_data_ins, lh_env_config))
            else if (lane_num == 3)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane3(lane_data_ins, lh_env_config))
            else if (lane_num == 4)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane4(lane_data_ins, lh_env_config))
            else if (lane_num == 5)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane5(lane_data_ins, lh_env_config))
            else if (lane_num == 6)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane6(lane_data_ins, lh_env_config))
            else if (lane_num == 7)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane7(lane_data_ins, lh_env_config))
            else if (lane_num == 8)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane8(lane_data_ins, lh_env_config))
            else if (lane_num == 9)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane9(lane_data_ins, lh_env_config))
            else if (lane_num == 10)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane10(lane_data_ins, lh_env_config))
            else if (lane_num == 11)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane11(lane_data_ins, lh_env_config))
            else if (lane_num == 12)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane12(lane_data_ins, lh_env_config))
            else if (lane_num == 13)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane13(lane_data_ins, lh_env_config))
            else if (lane_num == 14)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane14(lane_data_ins, lh_env_config))
            else if (lane_num == 15)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane15(lane_data_ins, lh_env_config))

          end //}

          tenb_8b_decode();

          // If IDLE2 is not truncated, 36 bytes after 4M of cs field
          // marker, the IDLE2 cs field will get completed. Hence, if another IDLE2
          // sequence starts with D0.0, it'll be properly descrambled.
	  // If this condition is executed at the end of the whole block, then cs field
	  // truncation at its last byte is not taken care. Because its idle2_cs will
	  // also be made '0', and the idle2_cs_field_descrambled_data would not be used
	  // in the rx_data_handler block. Moving the following logic here will take care
	  // of the issue, because idle2_cs will be cleared in the next posedge only.
          if (cs_field_byte_cnt == 36)
          begin //{
            lane_data_ins.idle2_cs = 0;
            cs_field_byte_cnt = 0;
          end //}
          if (lane_data_ins.character == SRIO_M && lane_data_ins.cntl)
          begin //{
            M_cnt++;
            if (M_cnt>1)
            begin
              lane_data_ins.idle2_cs = 1;
            end
          end //}
          else if (M_cnt>0)
            M_cnt = 0;

          // Once CS marker started, if either K or SC or PD is received, then it means CS field marker / cs field
          // is completed or truncated. IDLE2 marker or CS field check happens in IDLE2 checker in Rx data
          // handler class.
          if (lane_data_ins.idle2_cs == 1 && lane_data_ins.cntl && (lane_data_ins.character == SRIO_K || lane_data_ins.character == SRIO_SC || lane_data_ins.character == SRIO_PD))
          begin //{
            lane_data_ins.idle2_cs = 0;
            cs_field_byte_cnt = 0;
            if(lane_data_ins.cntl && (lane_data_ins.character == SRIO_K) &&  lh_trans.port_initialized)
             begin//{
              `uvm_error("SRIO_PL_LANE_HANDLER : IDLE2_CS_FIELD_TRUNCATED_WITH_K", $sformatf(" Spec reference 4.7.4. Lane number : %0d. Idle2 CS field is truncated with K", lane_num))
             end//}
          end //}
          else if (lane_data_ins.idle2_cs == 1 && ~lane_data_ins.cntl)
          begin //{

            cs_field_byte_cnt++; // counting only after 4M of cs field marker.

            if (cs_field_byte_cnt == 1 || cs_field_byte_cnt == 3)
            begin //{

              if (lane_data_ins.character !== SRIO_D21_5 && lane_data_ins.character !== SRIO_D10_2)
              begin //{

          	// IDLE2 truncated in CS marker.

                lane_data_ins.idle2_cs = 0;
                cs_field_byte_cnt = 0;

              end //}

            end //}
            else if (cs_field_byte_cnt > 4)
            begin //{

              // Checking Dx.y will add huge logic since there are lot of
              // combinations for it based on which mode it initialized and
              // which modes are supported etc. Hence, checking D21.5 and cs
              // field characters for truncation. It is good enough to detect
              // the idle2 truncation.


              // IDLE2 truncated in CS Field.

              if (lane_data_ins.character != 8'h67 && lane_data_ins.character != 8'h78 && lane_data_ins.character != 8'h7E && lane_data_ins.character != 8'hF8)
              begin //{
                lane_data_ins.idle2_cs = 0;
                cs_field_byte_cnt = 0;
              end //}

            end //}

          end //}

          //if (lh_env_config.srio_mode != SRIO_GEN13)
          //begin //{
          //  if (mon_type && ((lh_config.tx_scr_en && ~lh_trans.idle_detected) || (lh_config.tx_scr_en && lh_trans.idle_detected && lh_trans.idle_selected)))
          //    data_descramble();
          //  else if (~mon_type && ((lh_config.tx_scr_en && ~lh_trans.idle_detected) || (lh_config.tx_scr_en && lh_trans.idle_detected && lh_trans.idle_selected)))
          //    data_descramble();
          //end //}

          if (lh_env_config.srio_mode != SRIO_GEN13)
          begin //{

            if (mon_type && lh_env_config.srio_tx_mon_if == BFM)
            begin //{

              if ((lh_config.tx_scr_en && ~lh_trans.idle_detected) || (lh_config.tx_scr_en && lh_trans.idle_detected && lh_trans.idle_selected))
                data_descramble();

            end //}
            else if (mon_type && lh_env_config.srio_tx_mon_if == DUT)
            begin //{

	      register_update_method("Control_2_CSR", "Data_scrambling_disable", 64, "lh_reg_model_tx", reqd_field_name["Data_scrambling_disable"]);
	      dut_tx_scr_dis = reqd_field_name["Data_scrambling_disable"].get();
              //dut_tx_scr_dis = lh_env_config.srio_reg_model_tx.Port_0_Control_2_CSR.Data_scrambling_disable.get();
              if ((~dut_tx_scr_dis && ~lh_trans.idle_detected) || (~dut_tx_scr_dis && lh_trans.idle_detected && lh_trans.idle_selected))
                data_descramble();

            end //}

            if (~bfm_or_mon && ~mon_type && lh_env_config.srio_rx_mon_if == BFM)
            begin //{

              if ((lh_config.tx_scr_en && ~lh_trans.idle_detected) || (lh_config.tx_scr_en && lh_trans.idle_detected && lh_trans.idle_selected))
                data_descramble();

            end //}
            else if (~bfm_or_mon && ~mon_type && lh_env_config.srio_rx_mon_if == DUT)
            begin //{

	      register_update_method("Control_2_CSR", "Data_scrambling_disable", 64, "lh_reg_model_rx", reqd_field_name["Data_scrambling_disable"]);
	      dut_tx_scr_dis = reqd_field_name["Data_scrambling_disable"].get();
              //dut_tx_scr_dis = lh_env_config.srio_reg_model_rx.Port_0_Control_2_CSR.Data_scrambling_disable.get();
              if ((~dut_tx_scr_dis &&~lh_trans.idle_detected) || (~dut_tx_scr_dis && lh_trans.idle_detected && lh_trans.idle_selected))
                data_descramble();

            end //}

            if (bfm_or_mon)
            begin //{

              if ((lh_config.tx_scr_en && ~lh_trans.idle_detected) || (lh_config.tx_scr_en && lh_trans.idle_detected && lh_trans.idle_selected))
                data_descramble();

            end //}

          end //}



          //`uvm_info("SRIO_LANE_HANDLER : DESCRAMBLED DATA", $sformatf("LANE NUM : %0d Descrambled data is %0h", lane_num, lane_data_ins.character), UVM_LOW)

          if (lh_env_config.srio_interface_mode == SRIO_SERIAL)
            divide_clk = ~divide_clk;

        end //}

      end //}
      else
      begin //{  GEN3.0
	  if (lh_trans.frame_lock[lane_num])
	  begin //{
	    sixty_seven_bit_data = 67'h0_0000_0000_0000_0000;
            sixty_seven_bit_cnt = 0;
	    s2p_lock = 0;
            //divide_clk = 0;
            //note_bit_2=66;
            note_bit_1=67;
	  end //}

        if (lh_env_config.srio_interface_mode == SRIO_SERIAL)
        begin //{

          sixty_seven_bit_data = sixty_seven_bit_data<<1;
          sixty_seven_bit_data[66] = rx_data;

	  if (lh_trans.frame_lock[lane_num])
	  begin //{
	    sixty_seven_bit_data = 67'h0_0000_0000_0000_0000;
            sixty_seven_bit_cnt = 0;
	    s2p_lock = 0;
            divide_clk = 0;
	  end //}
	  else
            sixty_seven_bit_cnt++;

	  if (lh_config.brc3_training_mode)
	  begin //{
            dme_frame_sixty_seven_bit_data = dme_frame_sixty_seven_bit_data<<1;
            dme_frame_sixty_seven_bit_data[66] = rx_data;
	    dme_frame_sixty_seven_bit_cnt++;
		//$display($time, " dme_frame_sixty_seven_bit_cnt is %0d", dme_frame_sixty_seven_bit_cnt);
	  end //}

        end //}
        else if (lh_env_config.srio_interface_mode == SRIO_PARALLEL)
        begin //{

          if(~lh_config.parallel_cw_slip_adj_en || (!lh_trans.lane_trained[lane_num] && lh_config.brc3_training_mode))
           begin//{
          sixty_seven_bit_data = gen3_rx_pdata;
            if(~s2p_lock && ~lh_config.parallel_cw_slip_adj_en)
             begin//{
	        if (sixty_seven_bit_data[1] == ~sixty_seven_bit_data[2])
                 begin//{
	          s2p_lock = 1;
                 end//}
             end//}
           end//}
          else
           begin//{
          if(lh_env_config.srio_interface_mode == SRIO_PARALLEL && s2p_lock)
           begin//{
            sixty_seven_bit_data=sixty_seven_bit_data_tmp;
           end//}
            sixty_seven_bit_data_tmp = gen3_rx_pdata;
            if(~s2p_lock)
             begin//{
              for(int k=0;k<=note_bit_1;k++)
               begin//{
	        if (sixty_seven_bit_data[1] == ~sixty_seven_bit_data[2])
                 begin//{
	          s2p_lock = 1;
                  note_bit_1=k;
                  if(k==67)
                   note_bit_1=0;
//`uvm_info("LANE_HANDL",$sformatf("note_bit_1:%0d",note_bit_1),UVM_LOW)
                  break;
                 end//}
                else
                 begin//{
                  if(k!=67)
                   begin//{
                    sixty_seven_bit_data=sixty_seven_bit_data<<1;
                    sixty_seven_bit_data[66]=sixty_seven_bit_data_tmp[0];
                    sixty_seven_bit_data_tmp=sixty_seven_bit_data_tmp<<1;
//`uvm_info("LANE_HANDL",$sformatf("k:%0d sixty_seven_bit_data:%x,sixty_seven_bit_data_tmp:%x",k,sixty_seven_bit_data,sixty_seven_bit_data_tmp),UVM_LOW)
                   end//}
                 end//}
               end//}
            end//}
           else
            begin//{
              slice=67-note_bit_1;
              lsb=0;
              for(int i=slice;i<67;i++)
               begin//{
               sixty_seven_bit_data[i]=sixty_seven_bit_data_tmp[lsb];
               lsb++;
               end//}
              sixty_seven_bit_data_tmp=sixty_seven_bit_data_tmp<<note_bit_1;
            end//}
           end//}
//`uvm_info("LANE_HANDL",$sformatf(" sixty_seven_bit_data:%x,sixty_seven_bit_data_tmp:%x",sixty_seven_bit_data,sixty_seven_bit_data_tmp),UVM_LOW)

	  if (lh_config.brc3_training_mode)
           begin//{
             if(~lh_config.parallel_dme_slip_adj_en)
              dme_frame_sixty_seven_bit_data = gen3_rx_pdata;
             else
              begin//{
               dme_frame_sixty_seven_bit_data_tmp = gen3_rx_pdata;
               if(parallel_slide_mode)
                dme_frame_sixty_seven_bit_data = gen3_rx_pdata;
              end//}
           end//}
           if(lh_config.parallel_dme_slip_adj_en)
            gen3_rx_pdata=gen3_rx_pdata_tmp;

        end //}

        if (lh_env_config.srio_interface_mode == SRIO_SERIAL)
        begin //{

          if (sixty_seven_bit_cnt == 67 && ~s2p_lock)
          begin //{

	    if (sixty_seven_bit_data[1] == ~sixty_seven_bit_data[2])
	      s2p_lock = 1;
            else
              sixty_seven_bit_cnt--;

//          `uvm_info("SRIO_LANE_HANDLER :", $sformatf("LANE NUM : %0d 67 bit data is %0h", lane_num, sixty_seven_bit_data), UVM_LOW)

          end //}

	  
          if (dme_frame_sixty_seven_bit_cnt == 67 && ~dme_frame_s2p_lock)
          begin //{

	    if (lh_trans.dme_mode[lane_num] && dme_frame_sixty_seven_bit_data[0:31] == 32'hFFFF_0000) // Frame marker detection.
	      dme_frame_s2p_lock = 1;
            else
              dme_frame_sixty_seven_bit_cnt--;

	    if (dme_frame_s2p_lock)
	    begin //{

	      frame_marker_data = dme_frame_sixty_seven_bit_data[0:31];
	      new_marker = 1;

	    end //}

          end //}
	  else if (dme_frame_sixty_seven_bit_cnt == 67 && dme_frame_s2p_lock)
	  begin //{

	    if (current_frame_lock_state == SLIP)
	    begin //{
	      slip_done = 1;
	      frame_bit_count = 0;
	      frame_offset_achieved = 0;
	    end //}

	  end //}

          if (sixty_seven_bit_cnt == 33 && s2p_lock)
            divide_clk = ~divide_clk;

	  if (dme_frame_sixty_seven_bit_cnt == 33 && dme_frame_s2p_lock)
            dme_frame_divide_clk = ~dme_frame_divide_clk;

        end //}
	else
	begin //{

	  if (lh_config.brc3_training_mode && ~gen3_parallel_mode_frame_received)
	  begin //{
             if(~lh_config.parallel_dme_slip_adj_en)
              begin//{ 
	    if (dme_frame_sixty_seven_bit_data[0:31] == 32'hFFFF_0000)
	    begin //{

	      gen3_parallel_mode_frame_received = 1;
	      frame_marker_data = dme_frame_sixty_seven_bit_data[0:31];
	      new_marker = 1;

	    end //}
	   end //}
          else
	   begin //{
            for(int k=0;k<=(note_bit_2+1);k++)
             begin//{
              if(dme_frame_sixty_seven_bit_data[0:31] == 32'hFFFF_0000)
               begin//{
               note_bit_2=k;
               if(k==67)
                note_bit_2=0;
               gen3_rx_pdata=gen3_rx_pdata<<note_bit_2;
               break;
               end//}
              else
               begin//{
                if(k!=67)
                 begin//{
                  dme_frame_sixty_seven_bit_data=dme_frame_sixty_seven_bit_data<<1;
                  dme_frame_sixty_seven_bit_data[66]=dme_frame_sixty_seven_bit_data_tmp[0];
                  dme_frame_sixty_seven_bit_data_tmp=dme_frame_sixty_seven_bit_data_tmp<<1;
                 end//}
               end//}
             end//}
	    if (dme_frame_sixty_seven_bit_data[0:31] == 32'hFFFF_0000)
	    begin //{
              parallel_slide_mode=1;
	      gen3_parallel_mode_frame_received = 1;
	      frame_marker_data = dme_frame_sixty_seven_bit_data[0:31];
	      new_marker = 1;
	    end //}
	   end //}
          

	  end //}
	  else if (lh_config.brc3_training_mode && gen3_parallel_mode_frame_received)
	  begin //{

	    if (current_frame_lock_state == SLIP)
	    begin //{
	      slip_done = 1;
	      gen3_parallel_mode_frame_received = 0;
	      frame_bit_count = 0;
	      frame_offset_achieved = 0;
	    end //}

	  end //}

	end //}

        if ((dme_frame_sixty_seven_bit_cnt == 67 && dme_frame_s2p_lock) || (lh_env_config.srio_interface_mode == SRIO_PARALLEL && lh_config.brc3_training_mode && gen3_parallel_mode_frame_received))
        begin //{

          lh_trans.signal_detect[lane_num] = 1;

          if (lh_env_config.srio_interface_mode == SRIO_SERIAL)
            dme_frame_sixty_seven_bit_cnt = 0;

	  // When frame offset is achieved, there could be few bits left in the previous
	  // 67-bit frame data which belongs to the new frame. This assignment is done
	  // here before assigning the new sixty_seven_bit_data to the brc3_frame_data.
	  // Before overwriting the complete_dme_frame below with the new frame information,
	  // it should have been sampled by the long run training method.
	  if (frame_offset_achieved)
	  begin //{

	    temp_remaining_bits = remaining_bits_in_prev_frame;

	    for (int ndf=0; ndf<frame_bit_count; ndf++)
	    begin //{
	      complete_dme_frame[ndf] = brc3_frame_data[temp_remaining_bits];
	      temp_remaining_bits++;
	    end //}

	  end //}

          brc3_frame_data = dme_frame_sixty_seven_bit_data;

	  frame_bit_count = frame_bit_count + 67;

	  if (frame_bit_count >= 4384) // 4384 bits comprise the complete DME frame which is 548 octets.
	  begin //{

	    temp_frame_bit_count = frame_bit_count;
	    temp_frame_bit_count = temp_frame_bit_count - 4384;
	    remaining_bits_in_prev_frame = 67 - temp_frame_bit_count;
	    temp_remaining_bits = remaining_bits_in_prev_frame;

	    // Here part-select for complete_dme_frame and brc3_frame_data
	    // is completely variable dependent and it is not allowed by 
	    // the simulator. Thus, used the for-loop as work around here.
	    for (int rdf=0; rdf<remaining_bits_in_prev_frame; rdf++)
	    begin //{
	      complete_dme_frame[4384-temp_remaining_bits] = brc3_frame_data[rdf];
	      temp_remaining_bits--;
	    end //}

	    frame_offset = 1;
	    frame_offset_achieved = 1;

	    frame_bit_count = temp_frame_bit_count;

	  end //}
	  else
	  begin //{

	    complete_dme_frame[(frame_bit_count-67)+:67] = brc3_frame_data;

	    if (frame_offset_achieved)
	    begin //{

	      frame_offset_achieved = 0;

	      frame_marker_data = complete_dme_frame[0:31];
	      new_marker = 1;

	    end //}

	  end //}

          if (lh_env_config.srio_interface_mode == SRIO_SERIAL)
            dme_frame_divide_clk = ~dme_frame_divide_clk;

	end //}

        if ((sixty_seven_bit_cnt == 67 && s2p_lock) || (lh_env_config.srio_interface_mode == SRIO_PARALLEL && s2p_lock))
        begin //{

          lh_trans.signal_detect[lane_num] = 1;

          if (lh_env_config.srio_interface_mode == SRIO_SERIAL)
            sixty_seven_bit_cnt = 0;
          sixty_seven_bit_data_reg=sixty_seven_bit_data;
          if (sixty_seven_bit_data[0])
          begin //{
	    -> lh_trans.invert_bit_high;
	    sixty_seven_bit_data = ~sixty_seven_bit_data;
	    sixty_seven_bit_data[1] = ~sixty_seven_bit_data[1]; // Reverting back type and !type bits.
	    sixty_seven_bit_data[2] = ~sixty_seven_bit_data[2];
          end //}

  	  if (~bfm_or_mon && (sixty_seven_bit_data[1] == sixty_seven_bit_data[2]))
  	  begin //{
  	    update_error_detect_csr("DELIN_ERR");
  	  end //}

          lane_data_ins.brc3_cg = sixty_seven_bit_data;
          if(lh_env_config.srio_interface_mode == SRIO_PARALLEL && s2p_lock)
           begin//{
            sixty_seven_bit_data=sixty_seven_bit_data_reg;
           end//}

          if (bfm_or_mon)
          begin //{

            if (lane_num == 0)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane0(lane_data_ins, lh_env_config))
            else if (lane_num == 1)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane1(lane_data_ins, lh_env_config))
            else if (lane_num == 2)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane2(lane_data_ins, lh_env_config))
            else if (lane_num == 3)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane3(lane_data_ins, lh_env_config))
            else if (lane_num == 4)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane4(lane_data_ins, lh_env_config))
            else if (lane_num == 5)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane5(lane_data_ins, lh_env_config))
            else if (lane_num == 6)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane6(lane_data_ins, lh_env_config))
            else if (lane_num == 7)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane7(lane_data_ins, lh_env_config))
            else if (lane_num == 8)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane8(lane_data_ins, lh_env_config))
            else if (lane_num == 9)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane9(lane_data_ins, lh_env_config))
            else if (lane_num == 10)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane10(lane_data_ins, lh_env_config))
            else if (lane_num == 11)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane11(lane_data_ins, lh_env_config))
            else if (lane_num == 12)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane12(lane_data_ins, lh_env_config))
            else if (lane_num == 13)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane13(lane_data_ins, lh_env_config))
            else if (lane_num == 14)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane14(lane_data_ins, lh_env_config))
            else if (lane_num == 15)
              `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_cg_received_lane15(lane_data_ins, lh_env_config))

          end //}

          sixty_sevenb_sixty_fourb_decode();

          if (mon_type && lh_env_config.srio_tx_mon_if == BFM)
          begin //{

            if (lh_config.tx_scr_en)
              gen3_data_descramble();

          end //}
          else if (mon_type && lh_env_config.srio_tx_mon_if == DUT)
          begin //{

	    register_update_method("Control_2_CSR", "Data_scrambling_disable", 64, "lh_reg_model_tx", reqd_field_name["Data_scrambling_disable"]);
	    dut_tx_scr_dis = reqd_field_name["Data_scrambling_disable"].get();
            //dut_tx_scr_dis = lh_env_config.srio_reg_model_tx.Port_0_Control_2_CSR.Data_scrambling_disable.get();
            if (~dut_tx_scr_dis)
              gen3_data_descramble();

          end //}

          if (~bfm_or_mon && ~mon_type && lh_env_config.srio_rx_mon_if == BFM)
          begin //{

            if (lh_config.tx_scr_en)
              gen3_data_descramble();

          end //}
          else if (~bfm_or_mon && ~mon_type && lh_env_config.srio_rx_mon_if == DUT)
          begin //{

	    register_update_method("Control_2_CSR", "Data_scrambling_disable", 64, "lh_reg_model_rx", reqd_field_name["Data_scrambling_disable"]);
	    dut_tx_scr_dis = reqd_field_name["Data_scrambling_disable"].get();
            //dut_tx_scr_dis = lh_env_config.srio_reg_model_rx.Port_0_Control_2_CSR.Data_scrambling_disable.get();
            if (~dut_tx_scr_dis)
              gen3_data_descramble();

          end //}

          if (bfm_or_mon)
          begin //{

            if (lh_config.tx_scr_en)
              gen3_data_descramble();

          end //}


          //`uvm_info("SRIO_LANE_HANDLER : DESCRAMBLED DATA", $sformatf("LANE NUM : %0d Descrambled data is %0h", lane_num, lane_data_ins.character), UVM_LOW)

	  if (lh_trans.lane_sync[lane_num] && lane_data_ins.brc3_cntl_cw_type == DATA && ~trigger_os_check_methods)
	    trigger_os_check_methods = 1;
	  else if (~lh_trans.lane_sync[lane_num])
	    trigger_os_check_methods = 0;

	  if (trigger_os_check_methods)
	  begin //{

	    status_cntl_os_check_method();

	    descr_seed_os_check_method();

	    skip_os_check_method();

	  end //}

          if (lh_env_config.srio_interface_mode == SRIO_SERIAL)
            divide_clk = ~divide_clk;

        end //}

      end //}

    end //}

  end //}

endtask : ser2par


////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : tenb_8b_decode
/// Description : 10bit to 8bit decoder method. The 10bit data received is used to check if the
/// corresponding 8b data is available in the decoder array based on the current running disparity.
/// If the matching entry is not found, the codegroup is marked as invalid. If the invalid codegroup
/// count reaches 15, then the s2p_lock is cleared, so that 10bit lock has to happen from the start.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::tenb_8b_decode();

  int temp_10b_data;

  temp_10b_data = lane_data_ins.cg;

  if (lh_trans.data_pos_rd_array.exists(temp_10b_data) && lane_data_ins.curr_rd == POS)
  begin //{

    lane_data_ins.character = lh_trans.data_pos_rd_array[temp_10b_data];
    lane_data_ins.cntl = 0;
    lane_data_ins.invalid_cg = 0;
    calc_curr_rd(temp_10b_data);

    //`uvm_info("SRIO_LANE_HANDLER : 10B_8B INFO", $sformatf("LANE NUM : %0d 1st if of tenb_8b_decode. tenb_data is %0h 8b_char is %0h, CURRENT RUNNING DISPARITY is %0s", lane_num, temp_10b_data, lane_data_ins.character, lane_data_ins.curr_rd.name()), UVM_LOW)

    return;

  end //}

  if (lh_trans.data_neg_rd_array.exists(temp_10b_data) && lane_data_ins.curr_rd == NEG)
  begin //{

    lane_data_ins.character = lh_trans.data_neg_rd_array[temp_10b_data];
    lane_data_ins.cntl = 0;
    lane_data_ins.invalid_cg = 0;
    calc_curr_rd(temp_10b_data);

    //`uvm_info("SRIO_LANE_HANDLER :10B_8B INFO", $sformatf("LANE NUM : %0d 2nd if of tenb_8b_decode. tenb_data is %0h 8b_char is %0h, CURRENT RUNNING DISPARITY is %0s", lane_num, temp_10b_data, lane_data_ins.character, lane_data_ins.curr_rd.name()), UVM_LOW)

    return;

  end //}

  if (lh_trans.cntl_pos_rd_array.exists(temp_10b_data) && lane_data_ins.curr_rd == POS)
  begin //{

    lane_data_ins.character = lh_trans.cntl_pos_rd_array[temp_10b_data];
    lane_data_ins.cntl = 1;
    lane_data_ins.invalid_cg = 0;
    calc_curr_rd(temp_10b_data);

    //`uvm_info("SRIO_LANE_HANDLER :10B_8B INFO", $sformatf("LANE NUM : %0d 3rd if of tenb_8b_decode. tenb_data is %0h 8b_char is %0h, CURRENT RUNNING DISPARITY is %0s", lane_num, temp_10b_data, lane_data_ins.character, lane_data_ins.curr_rd.name()), UVM_LOW)

    return;

  end //}

  if (lh_trans.cntl_neg_rd_array.exists(temp_10b_data) && lane_data_ins.curr_rd == NEG)
  begin //{

    lane_data_ins.character = lh_trans.cntl_neg_rd_array[temp_10b_data];
    lane_data_ins.cntl = 1;
    lane_data_ins.invalid_cg = 0;
    calc_curr_rd(temp_10b_data);

    //`uvm_info("SRIO_LANE_HANDLER :10B_8B INFO", $sformatf("LANE NUM : %0d 4th if of tenb_8b_decode. tenb_data is %0h 8b_char is %0h, CURRENT RUNNING DISPARITY is %0s", lane_num, temp_10b_data, lane_data_ins.character, lane_data_ins.curr_rd.name()), UVM_LOW)

    return;

  end //}

  lane_data_ins.invalid_cg = 1;

// TODO:temp logic. clearing of s2p_lock logic has to be finalized. Also check if this logic itself holds good.
  invalid_cg_cnt++;

  if (invalid_cg_cnt == 15)
  begin //{
    s2p_lock = 0;
    invalid_cg_cnt = 0;
  end //}

  if (~bfm_or_mon)
  begin //{
    update_error_detect_csr("INVALID_CHAR");
  end //}

    //if (~bfm_or_mon && mon_type && lh_trans.port_initialized)
    //  `uvm_info("SRIO_LANE_HANDLER :10B_8B INFO", $sformatf("LANE NUM : %0d Invalid CG detected in tenb_8b_decode. tenb_data is %0h CURRENT RUNNING DISPARITY is %0s", lane_num, temp_10b_data, lane_data_ins.curr_rd.name()), UVM_LOW)

endtask : tenb_8b_decode


////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : calc_curr_rd
/// Description : Calculates the current running disparity. Logic follows the algorithm described in
/// section 4.5.3 of RIO2.2, Part6 specification.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::calc_curr_rd(input int data);

  bit [0:9] temp_data;

  bit left_part_ones_greater;
  bit right_part_ones_greater;

  bit ones_zeros_equal;

  int ones_cnt;
  int zeros_cnt;

  running_disparity curr_disp;

  ones_cnt = 0;
  zeros_cnt = 0;

  curr_disp = lane_data_ins.curr_rd;
  temp_data = data;

  for (int find_ones_cnt=0; find_ones_cnt<6; find_ones_cnt++)
  begin //{
    if (temp_data[find_ones_cnt] == 1)
      ones_cnt++;
    else
      zeros_cnt++;
  end //}

  if (ones_cnt > zeros_cnt)
    left_part_ones_greater = 1;
  else if (ones_cnt == zeros_cnt)
    ones_zeros_equal = 1;
  else 
    left_part_ones_greater = 0;


  if (left_part_ones_greater || (temp_data[0:5] == 6'b000111))
    curr_disp = POS;
  else if ((~left_part_ones_greater && ~ones_zeros_equal) || (temp_data[0:5] == 6'b111000))
    curr_disp = NEG;
  else
    curr_disp = curr_disp;

  ones_cnt = 0;
  zeros_cnt = 0;
  ones_zeros_equal = 0;

  for (int find_ones_cnt=6; find_ones_cnt<10; find_ones_cnt++)
  begin //{
    if (temp_data[find_ones_cnt] == 1)
      ones_cnt++;
    else
      zeros_cnt++;
  end //}

  if (ones_cnt > zeros_cnt)
    right_part_ones_greater = 1;
  else if (ones_cnt == zeros_cnt)
    ones_zeros_equal = 1;
  else
    right_part_ones_greater = 0;


  if (right_part_ones_greater || (temp_data[6:9] == 4'b0011))
    curr_disp = POS;
  else if ((~right_part_ones_greater && ~ones_zeros_equal) || (temp_data[6:9] == 4'b1100))
    curr_disp = NEG;
  else
    curr_disp = curr_disp;

  lane_data_ins.curr_rd = curr_disp;

endtask : calc_curr_rd


////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : data_descramble
/// Description : Descrambler method, used for GEN2.x. Method returns immediately if IDLE1 is
/// detected, or if SKIP character (R) is received as part of IDLE2 sequence. MDDDD sequence is used
/// to initialize the descrsambler lfsr and then everytime a 'M' character is received, this method
/// performs the descrambler sync check. Descrambler sync check is performed by checking that 4
/// consecutive 'D' characters following the 'M' character are descrambled to '0' or not. If the
/// sync check fails, then the descrambler lfsr is initialized again using the next MDDDD sequence.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::data_descramble();

    //`uvm_info("SRIO_LANE_HANDLER : DESCRAMBLER DEBUG", $sformatf("LANE NUM : %0d Start of data_descramble task. descr_in_sync is %0d, start_descr_sync is %0d, descr_sync_check is %0d idle2_cs is %0d, prev_idle2_cs is %0d. character & cntl is %0h %0d", lane_num, descr_in_sync, start_descr_sync, descr_sync_check, lane_data_ins.idle2_cs, prev_idle2_cs, lane_data_ins.character, lane_data_ins.cntl), UVM_LOW)

  if (lh_trans.idle_detected && ~lh_trans.idle_selected) // IDLE1 selected. Descrambling is skipped.
    return;

  if (lane_data_ins.character == SRIO_R && lane_data_ins.cntl) // Skip character received. Don't shift the lfsr
    return;

  // Initially wait for an 'M' character to be received, and then
  // start the descrambler sync process.
  if (~descr_in_sync && ~start_descr_sync && ~descr_sync_check)
  begin //{
    descr_lfsr = 17'h1_ffff;
    if (lane_data_ins.character == SRIO_M && lane_data_ins.cntl)
      start_descr_sync = 1;
    return;
  end //}

  // Once descrambler sync process is started, the 4 consecutive 'D'
  // characters are expected to initialize the descrambler LFSR, but
  // the received 'M' was a part of IDLE2 CS Marker field, then the
  // descrambler sync process should be dropped and wait for next 'M'
  // character to start the descrambler sync process again.
  if (start_descr_sync && lane_data_ins.idle2_cs && ~descr_in_sync)
  begin //{

    start_descr_sync = 0;
    return;

  end //}

  // Once the descrambler sync process is started, the next 4 characters
  // after an 'M' will be D0.0. When D0.0 is scrambled, it'll result in 
  // the LFSR value. Hence, 3 'D' characters are used to load the descrambler
  // LFSR, and then it is shifted 3 times, so that the 4th 'D' character, is 
  // descrambled to '0'. This is done in init_lfsr task. If the 4th 'D' character
  // is not '0', then descrambler sync process is repeated again. On the other hand, if
  // the 4th 'D' character is successfully descrambled to '0', then descrambler sync check
  // process is triggered.
  if (start_descr_sync && ~lane_data_ins.idle2_cs && ~descr_sync_check && ~lane_data_ins.cntl)
  begin //{
    D_after_M_cnt++;
    init_lfsr();
    lane_data_ins.character = descr_lfsr[16:9] ^ lane_data_ins.character; // data descrambling logic.

    if (D_after_M_cnt == 4)
    begin //{

      D_after_M_cnt = 0;

      if (lane_data_ins.character == SRIO_D00)
      begin //{

	start_descr_sync = 0;
	descr_sync_check = 1;

      end //}
      else
      begin //{
	start_descr_sync = 0;
      end //}

    end //}

  end //}
  else if (~start_descr_sync && descr_sync_check)
  begin //{

    if (lane_data_ins.cntl && lane_data_ins.character == SRIO_M && D_after_M_cnt == 0)
    begin //{
      shift_descr_lfsr();
      D_after_M_cnt++;
    end //}
    else if (D_after_M_cnt>0 && ~lane_data_ins.cntl && ~lane_data_ins.idle2_cs)
    begin //{

      // In descrambler sync check process, it is checked that the 4 'D' characters after
      // an 'M' character is successfully descrambled to '0' or not. 
      // If the descrambler sync check process successfully passes for 2 consecutive times,
      // then the descrambler is declared to be in sync, else, the descrambler sync process
      // is performed again.

      shift_descr_lfsr();
      lane_data_ins.character = descr_lfsr[16:9] ^ lane_data_ins.character; // data descrambling logic.
      D_after_M_cnt++;

      if (lane_data_ins.character != SRIO_D00)
      begin //{
	descr_sync_check = 0;
	D_after_M_cnt = 0;
      end //}
      else if (D_after_M_cnt == 5)
      begin //{
	D_after_M_cnt = 0;
	descr_sync_check_cnt++;
      end //}

      if (descr_sync_check_cnt == 2)
      begin //{
	descr_sync_check_cnt = 0;
	descr_sync_check = 0;
	descr_in_sync = 1;
      end //}

    end //}
    else
    begin //{

      shift_descr_lfsr();

      if (~lane_data_ins.cntl && ~lane_data_ins.idle2_cs)
        lane_data_ins.character = descr_lfsr[16:9] ^ lane_data_ins.character; // data descrambling logic.
      else if (~lane_data_ins.cntl && lane_data_ins.idle2_cs)
        lane_data_ins.idle2_cs_field_descrambled_data = descr_lfsr[16:9] ^ lane_data_ins.character; // data descrambling logic.

      if (D_after_M_cnt>0)
	D_after_M_cnt = 0; // clear it incase the above elseif condition had incremented it.

    end //}

  end //}
  else if (descr_in_sync)
  begin //{

    // Even when the descrambler is in sync, the sync check
    // is performed everytime an 'M' character is received,
    // which is not part of an IDLE2 CS field marker.

    shift_descr_lfsr();

    if (~lane_data_ins.cntl && ~lane_data_ins.idle2_cs)
      lane_data_ins.character = descr_lfsr[16:9] ^ lane_data_ins.character; // data descrambling logic.
    else if (~lane_data_ins.cntl && lane_data_ins.idle2_cs)
      lane_data_ins.idle2_cs_field_descrambled_data = descr_lfsr[16:9] ^ lane_data_ins.character; // data descrambling logic.

    if (lane_data_ins.cntl && lane_data_ins.character == SRIO_M && D_after_M_cnt == 0)
    begin //{
      D_after_M_cnt++;
    end //}
    else if (D_after_M_cnt>0 && ~lane_data_ins.cntl && lane_data_ins.idle2_cs)
    begin //{
      D_after_M_cnt = 0;
    end //}
    else if (D_after_M_cnt>0 && ~lane_data_ins.idle2_cs && prev_idle2_cs)
    begin //{
      // prev_idle2_cs will detect the idle2 truncation at cs marker or cs field level.
      // This logic will take care if cs marker is truncated right after 4Ms.
      D_after_M_cnt = 0;
    end //}
    else if (D_after_M_cnt>0 && ~lane_data_ins.cntl && ~lane_data_ins.idle2_cs && ~prev_idle2_cs)
    begin //{

      D_after_M_cnt++;

      if (lane_data_ins.character != SRIO_D00)
      begin //{
	descr_in_sync = 0;
	D_after_M_cnt = 0;

        if (~lh_trans.ies_state && lh_trans.link_initialized)
        begin //{
          lh_trans.ies_state = 1;
          lh_trans.ies_cause_value = 7;
	//$display($time, " 10. Vaidhy : ies_state set here");
        end //}

  	if (~bfm_or_mon)
  	begin //{
  	  update_error_detect_csr("DESCR_SYNC_LOSS");
  	end //}

      end //}
      else if (D_after_M_cnt == 5)
      begin //{
	D_after_M_cnt = 0;
      end //}

    end //}

  end //}
  prev_idle2_cs = lane_data_ins.idle2_cs;

endtask : data_descramble



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : init_lfsr
/// Description : It initializes the GEN2.x descrambler lfsr using the received MDDDD sequence.
/// data_descramble method will call this method when it receives the MDDDD sequence.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::init_lfsr();

  if (D_after_M_cnt == 1)
    descr_lfsr[16:9] = lane_data_ins.character;
  else if (D_after_M_cnt == 2)
    descr_lfsr[8:1] = lane_data_ins.character;
  else if (D_after_M_cnt == 3)
    descr_lfsr[0] = lane_data_ins.character[0];
  else if (D_after_M_cnt == 4)
  begin //{
    repeat(3)
      shift_descr_lfsr();
  end //}

endtask : init_lfsr



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : shift_descr_lfsr 
/// Description : When called, it shifts the GEN2.x descrambler lfsr by 8 times.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::shift_descr_lfsr();

  bit [7:0] temp_lfsr_byte;
  int temp_lfsr_byte_var;

  temp_lfsr_byte_var = 7;

  for (int lfsr_loop_var = 16; lfsr_loop_var >= 9; lfsr_loop_var--)
  begin //{
    temp_lfsr_byte[temp_lfsr_byte_var] = descr_lfsr[lfsr_loop_var] ^ descr_lfsr[lfsr_loop_var-9];
    temp_lfsr_byte_var--;
  end //}

  descr_lfsr = descr_lfsr<<8;
  descr_lfsr[7:0] = temp_lfsr_byte;

endtask : shift_descr_lfsr



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : lane_sync_sm
/// Description : Implements the lane_sync state machine for GEN13 and GEN2.x as per the respective
/// protocol. Waiting for the next negedge of clk or reset is bypassed when intermediate states are
/// encountered by the state machine.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::lane_sync_sm();

  //int K_counter;
  //int V_counter;
  //int I_counter;

#1;

  if (~srio_if.srio_rst_n)
  begin //{
    current_sync_state = NO_SYNC;
    if (~bfm_or_mon)
      current_sync_state_q.push_back(current_sync_state);
    // questasim and vcs doesn't work properly on associatuve array methods
    // Hence, a work-around is done here by setting the array values to 1 and
    // then clearing it immediately.
    lh_trans.lane_sync[lane_num] = 1;
    lh_trans.lane_sync[lane_num] = 0;

    lh_trans.rcvr_trained[lane_num] = 1;
    if (lh_config.aet_en)
      lh_trans.rcvr_trained[lane_num] = 0;

    lh_trans.signal_detect[lane_num] = 1;
    lh_trans.signal_detect[lane_num] = 0;
    lh_trans.lane_ready[lane_num] = 1;
    lh_trans.lane_ready[lane_num] = 0;
    lh_trans.from_sc_lane_ready[lane_num] = 1;
    lh_trans.from_sc_lane_ready[lane_num] = 0;
    K_counter = 0;
    V_counter = 0;
    I_counter = 0;
  end //}

  if (~bfm_or_mon)
    update_ls0_lane_num_field();

  forever
  begin //{

    // In the following conditions, there's no need to wait for the negedge of clock, 
    // as it would lead to missing of alternate data
    if (!(prev_sync_state == NO_SYNC_1 && current_sync_state == NO_SYNC_2) && !(prev_sync_state == NO_SYNC_3 && current_sync_state == NO_SYNC_2) && !(prev_sync_state == SYNC_1 && current_sync_state == SYNC_2) && !(prev_sync_state == SYNC_3 && current_sync_state == SYNC_2) && !(prev_sync_state == SYNC_4 && current_sync_state == SYNC_2))
      @(negedge divide_clk or negedge srio_if.srio_rst_n or negedge lh_trans.signal_detect[lane_num]);

    if (lh_trans.current_init_state == SILENT)
    begin //{
      parallel_slide_mode=0;
      current_sync_state = NO_SYNC;
      lh_trans.lane_sync[lane_num] = 0;
      K_counter = 0;
      V_counter = 0;
      I_counter = 0;
      note_bit_2=66;

      if (lh_config.aet_en)
        lh_trans.rcvr_trained[lane_num] = 0;

    end //}

    if (~srio_if.srio_rst_n || ~lh_trans.signal_detect[lane_num])
    begin //{

      prev_sync_state = current_sync_state;

      current_sync_state = NO_SYNC;

      lh_trans.lane_sync[lane_num] = 0;
      K_counter = 0;
      V_counter = 0;
      I_counter = 0;
      s2p_lock = 0;

      if (lh_config.aet_en)
        lh_trans.rcvr_trained[lane_num] = 0;

      if (~bfm_or_mon && prev_sync_state != current_sync_state)
	current_sync_state_q.push_back(current_sync_state);

    end //}
    else
    begin //{

      //`uvm_info("SRIO_LANE_HANDLER : SYNC_SM", $sformatf(" lane_sync[%0d] is %0d Present sync state is %0s", lane_num, lh_trans.lane_sync[lane_num], current_sync_state.name()), UVM_LOW)

      prev_sync_state = current_sync_state;

      case (current_sync_state)

	NO_SYNC : begin //{

		   //$display($time, " : Entered NO_SYNC in lane_num %0d", lane_num);

		     lh_trans.lane_sync[lane_num] = 0;
      		     K_counter = 0;
      		     V_counter = 0;
      		     I_counter = 0;

		     if (lh_env_config.srio_mode == SRIO_GEN13)
		     begin //{
		       if (lh_trans.signal_detect[lane_num] && `GEN1_COMMA_CHAR)
		         current_sync_state = NO_SYNC_1;
		     end //}
		     else
		     begin //{
		       if (lh_trans.signal_detect[lane_num] && `GEN2_COMMA_CHAR)
		         current_sync_state = NO_SYNC_1;
		     end //}

		   end //}

	NO_SYNC_1 : begin //{

		      lh_trans.lane_sync[lane_num] = 0;
      		      K_counter++;
      		      V_counter++;

		      if (lh_env_config.srio_mode == SRIO_GEN13)
		      begin //{

		        if (K_counter < lh_config.comma_cnt_threshold)
		          current_sync_state = NO_SYNC_2;
		        else if (K_counter == lh_config.comma_cnt_threshold)
		          current_sync_state = SYNC;

		      end //}
		      else
		      begin //{

		        if (K_counter < lh_config.comma_cnt_threshold || V_counter < lh_config.vmin_sync_threshold)
		          current_sync_state = NO_SYNC_2;
		        else if (K_counter > (lh_config.comma_cnt_threshold-1) && V_counter > (lh_config.vmin_sync_threshold-1))
		          current_sync_state = SYNC;

		      end //}

		    end //}

	NO_SYNC_2 : begin //{

		      lh_trans.lane_sync[lane_num] = 0;

		      if (lh_env_config.srio_mode == SRIO_GEN13)
		      begin //{

		        if (!`GEN1_COMMA_CHAR && ~lane_data_ins.invalid_cg)
		          current_sync_state = NO_SYNC_2;
		        else if (`GEN1_COMMA_CHAR && ~lane_data_ins.invalid_cg)
		          current_sync_state = NO_SYNC_1;
		        else if (lane_data_ins.invalid_cg)
		          current_sync_state = NO_SYNC;

		      end //}
		      else
		      begin //{

		        if (!`GEN2_COMMA_CHAR && ~lane_data_ins.invalid_cg)
		          current_sync_state = NO_SYNC_3;
		        else if (`GEN2_COMMA_CHAR && ~lane_data_ins.invalid_cg)
		          current_sync_state = NO_SYNC_1;
		        else if (lane_data_ins.invalid_cg)
		          current_sync_state = NO_SYNC;

		      end //}

		    end //}

	NO_SYNC_3 : begin //{

		      lh_trans.lane_sync[lane_num] = 0;
      		      V_counter++;

		      current_sync_state = NO_SYNC_2;

		    end //}

	SYNC : begin //{

	         lh_trans.lane_sync[lane_num] = 1;
      	         I_counter = 0;

		 if (~lane_data_ins.invalid_cg)
	           current_sync_state = SYNC;
		 else
	           current_sync_state = SYNC_1;

	       end //}

	SYNC_1 : begin //{

		   //$display($time, " : Entered SYNC_1 in lane_num %0d", lane_num);

	           lh_trans.lane_sync[lane_num] = 1;
      	           V_counter = 0;
      	           I_counter++;

		   if (I_counter < lh_config.sync_break_threshold)
	             current_sync_state = SYNC_2;
		   else
	             current_sync_state = NO_SYNC;

	       	 end //}

	SYNC_2 : begin //{

		   //$display($time, " : Entered SYNC_2 in lane_num %0d", lane_num);

	           lh_trans.lane_sync[lane_num] = 1;

		   if (~lane_data_ins.invalid_cg)
	             current_sync_state = SYNC_3;
		   else
	             current_sync_state = SYNC_1;

	       	 end //}

	SYNC_3 : begin //{

		   //$display($time, " : Entered SYNC_3 in lane_num %0d", lane_num);

	           lh_trans.lane_sync[lane_num] = 1;
      	           V_counter++;

		   if (V_counter < lh_config.valid_sync_threshold)
	             current_sync_state = SYNC_2;
		   else
	             current_sync_state = SYNC_4;

	       	 end //}

	SYNC_4 : begin //{

		   //$display($time, " : Entered SYNC_4 in lane_num %0d", lane_num);

	           lh_trans.lane_sync[lane_num] = 1;
      	           V_counter = 0;
      	           I_counter--;

		   if (I_counter > 0)
	             current_sync_state = SYNC_2;
		   else
	             current_sync_state = SYNC;

	       	 end //}

      endcase

      if (prev_sync_state != current_sync_state && (current_sync_state == SYNC || prev_sync_state == SYNC))
        `uvm_info("SRIO_LANE_HANDLER : SYNC_SM", $sformatf(" lane_sync[%0d] is %0d Next sync state is %0s", lane_num, lh_trans.lane_sync[lane_num], current_sync_state.name()), UVM_LOW)

      if (~bfm_or_mon && prev_sync_state != current_sync_state)
	current_sync_state_q.push_back(current_sync_state);

    end //}

    if (lh_trans.lane_sync[lane_num] == 1)
      begin
       temp_lane_data_ins = new lane_data_ins;
       //$cast(temp_lane_data_ins, lane_data_ins.clone());
       srio_rx_lane_event.trigger(temp_lane_data_ins);
      end
//	if (~bfm_or_mon && ~mon_type)
//	$display($time, " lane_num is %0d, mon_type is %0d. Event triggered from sync sm. lane_data_ins.character is %0h temp_lane_data_ins.character is %0h", lane_num, mon_type, lane_data_ins.character, temp_lane_data_ins.character);

  end //}

endtask : lane_sync_sm



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : lane_ready_gen
/// Description : Sets or clears the lane_ready signal for the available lanes based on the lane's
/// characteristics / capability to exchange data. Expressions used to set/clear lane_ready signal
/// is done based on the configured mode (SRIO_GEN13 / SRIO_GEN2.x / SRIO_GEN30). The value of lane
/// specific signals are stored in the common component transaction instance, so that it could be
/// used by any of the other components that has access to this common transaction instance. lane_ready
/// signal is used by the align and initialize state machines to settle in appropriate working mode.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::lane_ready_gen();

  wait(lh_trans.lane_sync.exists(lane_num) && lh_trans.rcvr_trained.exists(lane_num));

  forever begin //{

    if (lh_env_config.srio_mode != SRIO_GEN30)
    begin //{

      @(lh_trans.lane_sync[lane_num] or lh_trans.rcvr_trained[lane_num]);

      lh_trans.lane_ready[lane_num] = lh_trans.lane_sync[lane_num] & lh_trans.rcvr_trained[lane_num];

    end //}
    else
    begin //{

      @(lh_trans.lane_sync[lane_num] or lh_trans.lane_trained[lane_num] or lh_trans.lane_retraining[lane_num]);

      lh_trans.lane_ready[lane_num] = lh_trans.lane_sync[lane_num] & lh_trans.lane_trained[lane_num] & !lh_trans.lane_retraining[lane_num];
      lh_trans.from_sc_lane_ready[lane_num] = lh_trans.lane_ready[lane_num]; // TODO: temp assignment. Need to assign it from receiving status_cntl cw.

      //`uvm_info("LANE_READY DISPLAY", $sformatf(" lane_ready is %0d, lane_sync is %0d, lane_trained is %0d, lane_retraining is %0d", lh_trans.lane_ready[lane_num], lh_trans.lane_sync[lane_num], lh_trans.lane_trained[lane_num], lh_trans.lane_retraining[lane_num]), UVM_LOW)

    end //}

    if (~bfm_or_mon)
      update_other_ls0_fields();

  end //}

endtask : lane_ready_gen



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : collect_idle2_csfield
/// Description : Collects the IDLE2 CS field to perform adaptive equalization training and related
/// checks. The method runs forever, checks each character and detects the reception of CS field.
/// Once CS field is received, it decodes the CS field bytes into corresponding 2-bit data and pushes
/// it into cs_fld_char_q which will be process by the aet method. Once a complete CS field is received,
/// it also gives a hook for the srio_pl_aet_cs_received_lane<x> callbacks, so that the user can
/// modify the received CS field based on the test requirement.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::collect_idle2_csfield();

  if (~lh_config.aet_en)
    return;

  forever begin //{

    wait(lh_trans.idle_detected == 1 && lh_trans.idle_selected == 1 && lh_trans.rcvr_trained[lane_num] == 0);

    @(negedge divide_clk);

    if(lane_data_ins.character == SRIO_M && idle2_cs_fld_method_char_cnt == 0 && ~idle2_cs_field_started)
      idle2_cs_fld_method_char_cnt++;
    else if(lane_data_ins.character == SRIO_M && idle2_cs_fld_method_char_cnt == 1 && ~idle2_cs_field_started)
      idle2_cs_fld_method_char_cnt++;
    else if(lane_data_ins.character != SRIO_M && idle2_cs_fld_method_char_cnt == 1 && ~idle2_cs_field_started)
      idle2_cs_fld_method_char_cnt=0;
    else if(idle2_cs_fld_method_char_cnt > 1 && idle2_cs_fld_method_char_cnt < 8 && ~idle2_cs_field_started)
    begin //{
      idle2_cs_fld_method_char_cnt++;
      if (idle2_cs_fld_method_char_cnt == 6)
      begin //{

	idle2_cs_marker_port_width = lane_data_ins.character[0:2];
	idle2_cs_marker_lane_number = lane_data_ins.character[4:7]; // bits 8-11 in status_1_csr

      end //}
    end //}
    else if(idle2_cs_fld_method_char_cnt == 8 && ~idle2_cs_field_started && !(lane_data_ins.character == 8'h67 || lane_data_ins.character == 8'h78 || lane_data_ins.character == 8'h7E || lane_data_ins.character == 8'hF8))
      idle2_cs_fld_method_char_cnt=0; // IDLE2 sequence might be truncated.
    else if(idle2_cs_fld_method_char_cnt == 8 && ~idle2_cs_field_started && (lane_data_ins.character == 8'h67 || lane_data_ins.character == 8'h78 || lane_data_ins.character == 8'h7E || lane_data_ins.character == 8'hF8))
    begin //{

      idle2_cs_fld_method_char_cnt=0;
      idle2_cs_field_started = 1;

      lane_cs_fld_data_ins = new();

      if(lane_data_ins.character == 8'h67)
        lane_cs_fld_data_ins.cs_fld_char_q.push_back(2'b00);
      else if(lane_data_ins.character == 8'h78)
        lane_cs_fld_data_ins.cs_fld_char_q.push_back(2'b01);
      else if(lane_data_ins.character == 8'h7E)
        lane_cs_fld_data_ins.cs_fld_char_q.push_back(2'b10);
      else if(lane_data_ins.character == 8'hF8)
        lane_cs_fld_data_ins.cs_fld_char_q.push_back(2'b11);

    end //}
    else if(idle2_cs_field_started && (lane_data_ins.character == 8'h67 || lane_data_ins.character == 8'h78 || lane_data_ins.character == 8'h7E || lane_data_ins.character == 8'hF8))
    begin //{

      if(lane_data_ins.character == 8'h67)
        lane_cs_fld_data_ins.cs_fld_char_q.push_back(2'b00);
      else if(lane_data_ins.character == 8'h78)
        lane_cs_fld_data_ins.cs_fld_char_q.push_back(2'b01);
      else if(lane_data_ins.character == 8'h7E)
        lane_cs_fld_data_ins.cs_fld_char_q.push_back(2'b10);
      else if(lane_data_ins.character == 8'hF8)
        lane_cs_fld_data_ins.cs_fld_char_q.push_back(2'b11);

      if(lane_cs_fld_data_ins.cs_fld_char_q.size() == 32)
      begin //{

        idle2_aet_method();

	if (bfm_or_mon)
	begin //{

	  if (lane_num == 0)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane0(lane_cs_fld_data_ins))
	  else if (lane_num == 1)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane1(lane_cs_fld_data_ins))
	  else if (lane_num == 2)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane2(lane_cs_fld_data_ins))
	  else if (lane_num == 3)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane3(lane_cs_fld_data_ins))
	  else if (lane_num == 4)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane4(lane_cs_fld_data_ins))
	  else if (lane_num == 5)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane5(lane_cs_fld_data_ins))
	  else if (lane_num == 6)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane6(lane_cs_fld_data_ins))
	  else if (lane_num == 7)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane7(lane_cs_fld_data_ins))
	  else if (lane_num == 8)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane8(lane_cs_fld_data_ins))
	  else if (lane_num == 9)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane9(lane_cs_fld_data_ins))
	  else if (lane_num == 10)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane10(lane_cs_fld_data_ins))
	  else if (lane_num == 11)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane11(lane_cs_fld_data_ins))
	  else if (lane_num == 12)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane12(lane_cs_fld_data_ins))
	  else if (lane_num == 13)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane13(lane_cs_fld_data_ins))
	  else if (lane_num == 14)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane14(lane_cs_fld_data_ins))
	  else if (lane_num == 15)
            `uvm_do_callbacks(srio_pl_lane_handler, srio_pl_callback, srio_pl_aet_cs_received_lane15(lane_cs_fld_data_ins))

	end //}

      end //}

    end //}
    else if(idle2_cs_field_started && !(lane_data_ins.character == 8'h67 || lane_data_ins.character == 8'h78 || lane_data_ins.character == 8'h7E || lane_data_ins.character == 8'hF8))
    begin //{
      idle2_cs_field_started = 0;
      lane_cs_fld_data_ins.cs_fld_char_q.delete();
    end //}
    
  end //}

endtask : collect_idle2_csfield




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : idle2_aet_method
/// Description : This method will decode the received CS field data into different CS field
/// informations like training commands, status, ack, nak, receiver_trained, scrambling enable.
/// The decoded informations are assigned to respective common transaction fields by the bfm instance,
/// so that the transmit path can take appropriate action based on the received training command or
/// status if required. The monitor instance will trigger the related AET checks.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::idle2_aet_method();

  lane_cs_fld_data_ins.decode_idle2_cs_field_bits();    

  if (lane_cs_fld_data_ins.idle2_cs_fld_decode_success)
  begin //{

    if (lane_cs_fld_data_ins.idle2_cs_fld_cmd)
    begin //{

      lh_trans.idle2_aet_command_set[lane_num] = 1;

      if (lane_cs_fld_data_ins.idle2_cs_fld_tap_minus1_cmd != 2'b00)
      begin //{
        lh_trans.idle2_aet_cs_fld_tap_minus1_cmd[lane_num] = 1;
        lh_trans.idle2_aet_cs_fld_tap_minus1_cmd_val[lane_num] = lane_cs_fld_data_ins.idle2_cs_fld_tap_minus1_cmd;
      end //}
      else if (lane_cs_fld_data_ins.idle2_cs_fld_tap_plus1_cmd != 2'b00)
      begin //{
        lh_trans.idle2_aet_cs_fld_tap_plus1_cmd[lane_num] = 1;
        lh_trans.idle2_aet_cs_fld_tap_plus1_cmd_val[lane_num] = lane_cs_fld_data_ins.idle2_cs_fld_tap_plus1_cmd;
      end //}
      else if (lane_cs_fld_data_ins.idle2_cs_fld_reset_emp)
      begin //{
        lh_trans.idle2_aet_cs_fld_reset_cmd[lane_num] = 1;
      end //}
      else if (lane_cs_fld_data_ins.idle2_cs_fld_preset_emp)
      begin //{
        lh_trans.idle2_aet_cs_fld_preset_cmd[lane_num] = 1;
      end //}

    end //}
    else
    begin //{

      lh_trans.idle2_aet_command_set[lane_num] = 0;

      lh_trans.idle2_aet_cs_fld_tap_minus1_cmd[lane_num] = 0;
      lh_trans.idle2_aet_cs_fld_tap_plus1_cmd[lane_num] = 0;
      lh_trans.idle2_aet_cs_fld_reset_cmd[lane_num] = 0;
      lh_trans.idle2_aet_cs_fld_preset_cmd[lane_num] = 0;

    end //}

    lh_trans.idle2_aet_cs_fld_rcvr_trained[lane_num] = lane_cs_fld_data_ins.idle2_cs_fld_rcvr_trained;
    lh_trans.idle2_aet_cs_fld_data_scr_en[lane_num] = lane_cs_fld_data_ins.idle2_cs_fld_data_scr_en;
    lh_trans.idle2_aet_cs_fld_ack[lane_num] = lane_cs_fld_data_ins.idle2_cs_fld_ack;
    lh_trans.idle2_aet_cs_fld_nack[lane_num] = lane_cs_fld_data_ins.idle2_cs_fld_nack;

    if (~bfm_or_mon)
    begin //{

      if (prev_lane_cs_fld_data_ins != null)
      begin //{

	prev_lane_cs_fld_data_ins.compare_aet_control_fields(lane_cs_fld_data_ins);

	if (~prev_lane_cs_fld_data_ins.aet_fld_compare)
	  idle2_value_changed = 1;
	else
	begin //{

	  idle2_value_changed = 0;

	  prev_lane_cs_fld_data_ins.compare_aet_status_fields(lane_cs_fld_data_ins);

	  if (~prev_lane_cs_fld_data_ins.aet_fld_compare)
	    idle2_value_changed = 1;
	  else
	    idle2_value_changed = 0;

	end //}

      end //}

      lane_status_1_reg_val = {15'h0000, lane_cs_fld_data_ins.idle2_cs_fld_data_scr_en, lane_cs_fld_data_ins.idle2_cs_fld_tap_plus1_status[1], lane_cs_fld_data_ins.idle2_cs_fld_tap_plus1_status[0], lane_cs_fld_data_ins.idle2_cs_fld_tap_minus1_status[1], lane_cs_fld_data_ins.idle2_cs_fld_tap_minus1_status[0], idle2_cs_marker_lane_number[3], idle2_cs_marker_lane_number[2], idle2_cs_marker_lane_number[1], idle2_cs_marker_lane_number[0], idle2_cs_marker_port_width[2], idle2_cs_marker_port_width[1], idle2_cs_marker_port_width[0], lane_cs_fld_data_ins.idle2_cs_fld_rcvr_trained, 1'b0, idle2_value_changed, 2'b11};

      update_ls1_reg();

      prev_lane_cs_fld_data_ins = new lane_cs_fld_data_ins;

    end //}

    if (~bfm_or_mon)
      idle2_aet_checks();

  end //}

endtask : idle2_aet_method




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : idle2_aet_checks
/// Description : This method will perform the IDLE2 AET checks.
/// This method is triggered only by the monitor instance. The checks listed in the micro architecture
/// document under the section "PL monitor checks" and "AET checks" sub-section are covered in this
/// method.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::idle2_aet_checks();

  if ((mon_type && lh_env_config.srio_tx_mon_if == BFM) || (~mon_type && lh_env_config.srio_rx_mon_if == BFM))
  begin //{

    if (~lh_config.aet_en && lane_cs_fld_data_ins.idle2_cs_fld_cmd)
    begin //{

      `uvm_error("SRIO_PL_LANE_HANDLER: AET_ENABLE_CHECK", $sformatf(" Spec reference 6.6.10 / Table 6-18. Lane number is %0d. AET not supported, but equalization command transmitted", lane_num))

    end //}

  end //}
  else if ((mon_type && lh_env_config.srio_tx_mon_if == DUT) || (~mon_type && lh_env_config.srio_rx_mon_if == DUT))
  begin //{

    if (mon_type && lh_env_config.srio_tx_mon_if == DUT)
    begin //{
      register_update_method("Control_2_CSR", "Remote_Transmit_Emphasis_Control_Support", 64, "lh_reg_model_tx", reqd_field_name["Remote_Transmit_Emphasis_Control_Support"]);
      dut_rcvr_trn_spt = reqd_field_name["Remote_Transmit_Emphasis_Control_Support"].get();
      //dut_rcvr_trn_spt = lh_env_config.srio_reg_model_tx.Port_0_Control_2_CSR.Remote_Transmit_Emphasis_Control_Support.get();
      register_update_method("Control_2_CSR", "Remote_Transmit_Emphasis_Control_Enable", 64, "lh_reg_model_tx", reqd_field_name["Remote_Transmit_Emphasis_Control_Enable"]);
      dut_rcvr_trn_en = reqd_field_name["Remote_Transmit_Emphasis_Control_Enable"].get();
      //dut_rcvr_trn_en = lh_env_config.srio_reg_model_tx.Port_0_Control_2_CSR.Remote_Transmit_Emphasis_Control_Enable.get();
    end //}
    else if (~mon_type && lh_env_config.srio_rx_mon_if == DUT)
    begin //{
      register_update_method("Control_2_CSR", "Remote_Transmit_Emphasis_Control_Support", 64, "lh_reg_model_rx", reqd_field_name["Remote_Transmit_Emphasis_Control_Support"]);
      dut_rcvr_trn_spt = reqd_field_name["Remote_Transmit_Emphasis_Control_Support"].get();
      //dut_rcvr_trn_spt = lh_env_config.srio_reg_model_rx.Port_0_Control_2_CSR.Remote_Transmit_Emphasis_Control_Support.get();
      register_update_method("Control_2_CSR", "Remote_Transmit_Emphasis_Control_Enable", 64, "lh_reg_model_rx", reqd_field_name["Remote_Transmit_Emphasis_Control_Enable"]);
      dut_rcvr_trn_en = reqd_field_name["Remote_Transmit_Emphasis_Control_Enable"].get();
      //dut_rcvr_trn_en = lh_env_config.srio_reg_model_rx.Port_0_Control_2_CSR.Remote_Transmit_Emphasis_Control_Enable.get();
    end //}

    if (!(dut_rcvr_trn_spt && dut_rcvr_trn_en) && lane_cs_fld_data_ins.idle2_cs_fld_cmd)
    begin //{

      `uvm_error("SRIO_PL_LANE_HANDLER: AET_ENABLE_CHECK", $sformatf(" Spec reference 6.6.10 / Table 6-18. Lane number is %0d. AET not supported, but equalization command transmitted", lane_num))

    end //}
      
  end //}

  if (lane_cs_fld_data_ins.idle2_cs_fld_cmd)
  begin //{

    idle2_aet_cmd_cnt = 0;

    if (lane_cs_fld_data_ins.idle2_cs_fld_tap_minus1_cmd != 2'b00)
      idle2_aet_cmd_cnt++;

    if (lane_cs_fld_data_ins.idle2_cs_fld_tap_plus1_cmd != 2'b00)
      idle2_aet_cmd_cnt++;

    if (lane_cs_fld_data_ins.idle2_cs_fld_reset_emp)
      idle2_aet_cmd_cnt++;

    if (lane_cs_fld_data_ins.idle2_cs_fld_preset_emp)
      idle2_aet_cmd_cnt++;

    if (idle2_aet_cmd_cnt > 1)
    begin //{

      `uvm_error("SRIO_PL_LANE_HANDLER: AET_MULTIPLE_CMD_CHECK", $sformatf(" Spec reference 4.7.4.1.4. Lane number is %0d. More than one command set in the IDLE2 CS FIELD. TAP(-1) command is %0h, TAP(+1) command is %0h, Reset emphasis is %0h, Preset emphasis is %0h", lane_num, lane_cs_fld_data_ins.idle2_cs_fld_tap_minus1_cmd, lane_cs_fld_data_ins.idle2_cs_fld_tap_plus1_cmd, lane_cs_fld_data_ins.idle2_cs_fld_reset_emp, lane_cs_fld_data_ins.idle2_cs_fld_preset_emp))

    end //}

    idle2_aet_cmd_cnt = 0;

  end //}

  if (lane_cs_fld_data_ins.idle2_cs_fld_ack && lane_cs_fld_data_ins.idle2_cs_fld_nack)
  begin //{

    `uvm_error("SRIO_PL_LANE_HANDLER: AET_ACK_NACK_SET_CHECK", $sformatf(" Spec reference 4.7.4.1.4. Lane number is %0d. ACK and NACK are set together in a single IDLE2 CS FIELD", lane_num))

  end //}


  if (lane_cs_fld_data_ins.idle2_cs_fld_cmd || lane_cs_fld_data_ins.idle2_cs_fld_ack || lane_cs_fld_data_ins.idle2_cs_fld_nack)
  begin //{

    if (lane_cs_fld_data_ins.idle2_cs_fld_ack || lane_cs_fld_data_ins.idle2_cs_fld_nack)
    begin //{

      // This check will also catch the scenario when ACK/NACK
      //  is not de-asserted even after AET ACK/NACK timeout.
      if (~lh_common_mon_trans.idle2_aet_cmd_outstanding[~mon_type][lane_num])
      begin //{

    	`uvm_error("SRIO_PL_LANE_HANDLER: AET_ACK_WITHOUT_CMD_CHECK", $sformatf(" Spec reference 4.7.4.1.4. Lane number is %0d. ACK / NACK is set in IDLE2 CS FIELD when no AET command is outstanding, ACK is %0h, NACK is %0h", lane_num, lane_cs_fld_data_ins.idle2_cs_fld_ack, lane_cs_fld_data_ins.idle2_cs_fld_nack))

      end //}
      else
      begin //{
	lh_common_mon_trans.idle2_aet_ack_nack_rcvd[mon_type][lane_num] = 1;
      end //}

    end //}
    else if (lh_common_mon_trans.idle2_aet_ack_nack_rcvd[~mon_type][lane_num])
    begin //{
	// This else if block will get executed when the inbound aet command
	// ack process gets completed and at the same time it issues an outbound
	// aet command to its link partner.
      lh_common_mon_trans.idle2_aet_ack_nack_rcvd[~mon_type][lane_num] = 0;
    end //}

    if (~lh_common_mon_trans.idle2_aet_cmd_outstanding[mon_type][lane_num])
    begin //{

      if (lane_cs_fld_data_ins.idle2_cs_fld_cmd)
      begin //{

	if (check_cmd_reassertion && ~cmd_reassertion_timer_done)
	begin //{

    	  `uvm_error("SRIO_PL_LANE_HANDLER: AET_CMD_REASSERTION_CHECK", $sformatf(" Spec reference 4.7.4.1.4. Lane number is %0d. AET Command re-asserted before cmd_reassertion_timer_done.", lane_num))

	end //}

        bkp_lane_cs_fld_data_ins = new lane_cs_fld_data_ins;
        lh_common_mon_trans.idle2_aet_cmd_outstanding[mon_type][lane_num]= 1;

      end //}

    end //}
    else
    begin //{

      if (lh_common_mon_trans.idle2_ack_timeout_occured[~mon_type][lane_num])
      begin //{
      
        bkp_lane_cs_fld_data_ins.idle2_cs_fld_cmd = 0;
      
      end //}

      if (bkp_lane_cs_fld_data_ins.idle2_cs_fld_cmd && ~lh_common_mon_trans.idle2_aet_ack_nack_rcvd[~mon_type][lane_num])
      begin //{

	bkp_lane_cs_fld_data_ins.compare_aet_control_fields(lane_cs_fld_data_ins);

	if(~bkp_lane_cs_fld_data_ins.aet_fld_compare)
	begin //{

    	  `uvm_error("SRIO_PL_LANE_HANDLER: AET_CMD_CHANGE_BEFORE_ACK_CHECK", $sformatf(" Spec reference 4.7.4.1.4. Lane number is %0d. IDLE2 CS field command shall not change when neither ACK/NACK received nor AET command timeout occured. Expected command is %0h, Received command is %0h.    Expected tap_minus1_cmd is %0h, Received tap_minus1_cmd is %0h.   Expected tap_plus1_cmd is %0h, Received tap_plus1_cmd is %0h.     Expected Reset emphasis field is %0h, Received Reset emphasis field is %0h.     Expected Preset emphasis field is %0h, Received Preset emphasis field is %0h", lane_num, bkp_lane_cs_fld_data_ins.idle2_cs_fld_cmd, lane_cs_fld_data_ins.idle2_cs_fld_cmd, bkp_lane_cs_fld_data_ins.idle2_cs_fld_tap_minus1_cmd, lane_cs_fld_data_ins.idle2_cs_fld_tap_minus1_cmd, bkp_lane_cs_fld_data_ins.idle2_cs_fld_tap_plus1_cmd, lane_cs_fld_data_ins.idle2_cs_fld_tap_plus1_cmd, bkp_lane_cs_fld_data_ins.idle2_cs_fld_reset_emp, lane_cs_fld_data_ins.idle2_cs_fld_reset_emp, bkp_lane_cs_fld_data_ins.idle2_cs_fld_preset_emp, lane_cs_fld_data_ins.idle2_cs_fld_preset_emp))

	end //}

      end //}
      else if (bkp_lane_cs_fld_data_ins.idle2_cs_fld_cmd && lh_common_mon_trans.idle2_aet_ack_nack_rcvd[~mon_type][lane_num])
      begin //{

	if (~lane_cs_fld_data_ins.idle2_cs_fld_cmd)
	begin //{
	  bkp_lane_cs_fld_data_ins.idle2_cs_fld_cmd = 0;
	  lh_common_mon_trans.command_deasserted[mon_type][lane_num] = 1;
	end //}
	else if (lh_common_mon_trans.idle2_cmd_timeout_occured[mon_type][lane_num])
	begin //{

	  bkp_lane_cs_fld_data_ins.idle2_cs_fld_cmd = 0;

    	  `uvm_error("SRIO_PL_LANE_HANDLER: AET_CMD_DEASSERTION_AFTER_CMD_TIMEOUT_CHECK", $sformatf(" Spec reference 4.7.4.1.4. Lane number is %0d. AET Command not de-asserted even after command timeout occured.", lane_num))

	end //}

      end //}
      else if (~bkp_lane_cs_fld_data_ins.idle2_cs_fld_cmd && lane_cs_fld_data_ins.idle2_cs_fld_cmd && lh_common_mon_trans.idle2_ack_timeout_occured[~mon_type][lane_num])
      begin //{

    	`uvm_error("SRIO_PL_LANE_HANDLER: AET_CMD_DEASSERTION_AFTER_ACK_TIMEOUT_CHECK", $sformatf(" Spec reference 4.7.4.1.4. Lane number is %0d. AET Command not de-asserted after ACK timeout occured.", lane_num))

      end //}

    end //}

  end //}
  else
  begin //{

    if (lh_common_mon_trans.idle2_aet_ack_nack_rcvd[~mon_type][lane_num])
    begin //{

      if (bkp_lane_cs_fld_data_ins.idle2_cs_fld_cmd && ~lane_cs_fld_data_ins.idle2_cs_fld_cmd)
      begin //{

	bkp_lane_cs_fld_data_ins.idle2_cs_fld_cmd = 0;
	lh_common_mon_trans.command_deasserted[mon_type][lane_num] = 1;

      end //}

      //lh_common_mon_trans.idle2_aet_ack_nack_rcvd[~mon_type][lane_num] = 0;

    end //}
    else if (lh_common_mon_trans.idle2_aet_cmd_outstanding[mon_type][lane_num] && ~lh_common_mon_trans.idle2_aet_ack_nack_rcvd[~mon_type][lane_num] && ~lh_common_mon_trans.idle2_ack_timeout_occured[~mon_type][lane_num])
    begin //{

      `uvm_error("SRIO_PL_LANE_HANDLER: AET_CMD_DEASSERTION_BEFORE_ACK_CHECK", $sformatf(" Spec reference 4.7.4.1.4. Lane number is %0d. AET Command de-asserted unexpectedly when neither ack/nack received nor ack timeout occured.", lane_num))

    end //}

  end //}

endtask : idle2_aet_checks



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : set_receiver_trained
/// Description : This method will set the receiver_trained signal for SRIO_GEN2.x and lane_trained
/// and lane_retraining signals for SRIO_GEN30. The logic will run a timer and if any training
/// command is received before the timer expires, the timer is reloaded to the initial value.
/// This logic is implemented based on the assumption that training commands will not be required 
/// to be exchanged anymore if the lane is trained properly. Thus, receiver_trained or lane_trained 
/// signals will be set, only if no commands are detected till the timer expires.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::set_receiver_trained();

  if (lh_env_config.srio_mode != SRIO_GEN30)
  begin //{

    if (~lh_config.aet_en)
      return;

    lh_trans.idle2_aet_command_set[lane_num] = 1;
    lh_trans.idle2_aet_command_set[lane_num] = 0;

  end //}

    lh_trans.idle2_bfm_aet_command_set[lane_num] = 1;
    lh_trans.idle2_bfm_aet_command_set[lane_num] = 0;

    lh_trans.gen3_bfm_training_command_set[lane_num] = 1;
    lh_trans.gen3_bfm_training_command_set[lane_num] = 0;

  forever begin //{

    if (lh_env_config.srio_mode != SRIO_GEN30)
    begin //{

      wait(lh_trans.lane_sync[lane_num] == 1);
      wait(lh_trans.idle_detected == 1 && lh_trans.idle_selected == 1);

    end //}
    else
    begin //{

      wait(lh_trans.lane_sync[lane_num] == 1 || lh_trans.frame_lock[lane_num] == 1);

    end //}

    `uvm_info(" SRIO_PL_LANE_HANDLER : RECEIVER TRAINED TIMER", $sformatf(" STARTED for lane no. %0d", lane_num), UVM_LOW)

    if (~bfm_or_mon)
    begin //{

      repeat(lh_config.aet_training_period)
      begin //{

	if (lh_env_config.srio_mode != SRIO_GEN30)
	begin //{

          if (~lh_trans.idle2_aet_command_set[lane_num])
            @(posedge srio_if.sim_clk);
          else
            break;

	end //}
	else
	begin //{

          if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
            @(posedge srio_if.sim_clk);
          else
            break;

	end //}

      end //}

      if (lh_env_config.srio_mode != SRIO_GEN30)
      begin //{

        if (~lh_trans.idle2_aet_command_set[lane_num])
        begin //{

          lh_trans.rcvr_trained[lane_num] = 1;

          `uvm_info(" SRIO_PL_LANE_HANDLER : RECEIVER TRAINED TIMER", $sformatf(" ENDED. Receiver trained for lane no. %0d set.", lane_num), UVM_LOW)

        end //}
        else
          wait(lh_trans.idle2_aet_command_set[lane_num] == 0);

      end //}
      else
      begin //{

	// If cmd is outstanding in tx_monitor, it means, BFM is
	// transmitting cmd to train its local receiver. Thus, rx_monitor's
	// lane_trained signal has to be modified based on it. This is
	// done by checking gen3_training_cmd_outstanding[~mon_type] below.
        if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
        begin //{

          lh_trans.lane_trained[lane_num] = 1;
          lh_trans.lane_retraining[lane_num] = 0;

      	  lh_trans.from_sc_lane_trained[lane_num] = lh_trans.lane_trained[lane_num]; // TODO: temp assignment. Need to assign it from receiving status_cntl cw.

          `uvm_info(" SRIO_PL_LANE_HANDLER : RECEIVER TRAINED TIMER", $sformatf(" ENDED. Receiver trained for lane no. %0d set.", lane_num), UVM_LOW)

        end //}
        else
	begin //{
          lh_trans.lane_retraining[lane_num] = (lh_trans.retrain_lane[lane_num]) ? 1 : 0;
          wait(lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num] == 0);
	end //}

      end //}

    end //}
    else if (bfm_or_mon)
    begin //{

 // TODO: Add condition for srio_mode == SRIO_GEN30 once the signal is added in the TX_path

      if (lh_env_config.srio_mode != SRIO_GEN30)
      begin //{

        repeat(lh_config.aet_training_period)
        begin //{
          if (~lh_trans.idle2_bfm_aet_command_set[lane_num])
            @(posedge srio_if.sim_clk);
          else
            break;
        end //}

      end //}
      else if (lh_env_config.srio_mode == SRIO_GEN30)
      begin //{

        repeat(lh_config.aet_training_period)
        begin //{
          if (~lh_trans.gen3_bfm_training_command_set[lane_num])
            @(posedge srio_if.sim_clk);
          else
            break;
        end //}

      end //}

      if (lh_env_config.srio_mode != SRIO_GEN30)
      begin //{

        if (~lh_trans.idle2_bfm_aet_command_set[lane_num])
        begin //{

          lh_trans.rcvr_trained[lane_num] = 1;

          `uvm_info(" SRIO_PL_LANE_HANDLER : RECEIVER TRAINED TIMER", $sformatf(" ENDED. Receiver trained for lane no. %0d set.", lane_num), UVM_LOW)

        end //}
        else
        begin //{

          wait(lh_trans.idle2_bfm_aet_command_set[lane_num] == 0);

        end //}

      end //}
      else if (lh_env_config.srio_mode == SRIO_GEN30)
      begin //{

        if (~lh_trans.gen3_bfm_training_command_set[lane_num])
        begin //{

          lh_trans.lane_trained[lane_num] = 1;
          lh_trans.from_sc_lane_trained[lane_num] = lh_trans.lane_trained[lane_num]; // TODO: temp assignment. Need to assign it from receiving status_cntl cw.
          lh_trans.lane_retraining[lane_num] = 0;

          `uvm_info(" SRIO_PL_LANE_HANDLER : RECEIVER TRAINED TIMER", $sformatf(" ENDED. Receiver trained for lane no. %0d set.", lane_num), UVM_LOW)

        end //}
        else
        begin //{

          lh_trans.lane_retraining[lane_num] = (lh_trans.retrain_lane[lane_num]) ? 1 : 0;

          wait(lh_trans.gen3_bfm_training_command_set[lane_num] == 0);

        end //}

      end //}

    end //}

    if (lh_env_config.srio_mode != SRIO_GEN30)
    begin //{

      if (lh_trans.rcvr_trained[lane_num] == 1)
        wait(lh_trans.rcvr_trained[lane_num] == 0);

    end //}
    else
    begin //{

      if (lh_trans.lane_trained[lane_num] == 1)
        wait(lh_trans.lane_trained[lane_num] == 0);

    end //}

  end //}

endtask : set_receiver_trained



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : idle2_aet_timer_method
/// Description : This method runs different timers based on the current status of AET, such as
/// ack/nack timeout timer, command deassertion timer, ack/nack deassertion timer and command
/// reassertion timer in case of ack/nack timeout.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::idle2_aet_timer_method();

  if (~lh_config.aet_en)
    return;

  fork

    begin //{  ACK/NACK timeout logic

      forever begin //{

	wait(lh_common_mon_trans.idle2_aet_cmd_outstanding[mon_type][lane_num] == 1);

	repeat(lh_config.cs_field_ack_timer)
	begin //{
	  if (~lh_common_mon_trans.idle2_aet_ack_nack_rcvd[~mon_type][lane_num])
	    @(posedge srio_if.sim_clk);
	  else
	    break;
	end //}

	if (~lh_common_mon_trans.idle2_aet_ack_nack_rcvd[~mon_type][lane_num])
	begin //{
	  lh_common_mon_trans.idle2_ack_timeout_occured[~mon_type][lane_num] = 1;
	  check_cmd_reassertion = 1;
	end //}
	else
	  check_cmd_deassertion = 1;

	wait(lh_common_mon_trans.idle2_aet_cmd_outstanding[mon_type][lane_num] == 0);

      end //}

    end //}

    begin //{  CMD timeout logic

      forever begin //{

	wait(check_cmd_deassertion == 1);

	repeat(lh_config.aet_command_period)
	begin //{
	  if (~lh_common_mon_trans.command_deasserted[mon_type][lane_num])
	    @(posedge srio_if.sim_clk);
	  else
	    break;
	end //}

	if (~lh_common_mon_trans.command_deasserted[mon_type][lane_num])
	  lh_common_mon_trans.idle2_cmd_timeout_occured[mon_type][lane_num] = 1;

	lh_common_mon_trans.command_deasserted[mon_type][lane_num] = 0;
	check_cmd_deassertion = 0;

      end //}

    end //}

    begin //{  ACK/NACK deassertion logic

      forever begin //{

	wait(lh_common_mon_trans.idle2_aet_ack_nack_rcvd[mon_type][lane_num] == 1);
	wait(lh_common_mon_trans.command_deasserted[~mon_type][lane_num] == 1);

	repeat(lh_config.cs_field_ack_timer)
	begin //{
	  if (lh_common_mon_trans.idle2_aet_ack_nack_rcvd[mon_type][lane_num])
	    @(posedge srio_if.sim_clk);
	  else
	    break;
	end //}

	if (lh_common_mon_trans.idle2_aet_ack_nack_rcvd[mon_type][lane_num])
	  lh_common_mon_trans.idle2_aet_ack_nack_rcvd[mon_type][lane_num] = 0;

	cmd_reassertion_timer_done = 0;

	lh_common_mon_trans.idle2_cmd_timeout_occured[~mon_type][lane_num] = 0;
	lh_common_mon_trans.idle2_ack_timeout_occured[mon_type][lane_num] = 0;
	lh_common_mon_trans.idle2_aet_cmd_outstanding[~mon_type][lane_num] = 0;

      end //}

    end //}

    begin //{  CMD reassertion logic

      forever begin //{

	wait(check_cmd_reassertion == 1);
	cmd_reassertion_timer_done = 0;

	repeat(lh_config.aet_command_period)
	begin //{
	    @(posedge srio_if.sim_clk);
	end //}

	check_cmd_reassertion = 0;
	cmd_reassertion_timer_done = 1;

      end //}

    end //}

  join

endtask : idle2_aet_timer_method




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_ls0_lane_num_field
/// Description : This method updates the lane number field in the LaneN_Status_0 CSR.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_ls0_lane_num_field();

  if (lane_num == 0)
    void'(lh_reg_model.Lane_0_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 1)
    void'(lh_reg_model.Lane_1_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 2)
    void'(lh_reg_model.Lane_2_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 3)
    void'(lh_reg_model.Lane_3_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 4)
    void'(lh_reg_model.Lane_4_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 5)
    void'(lh_reg_model.Lane_5_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 6)
    void'(lh_reg_model.Lane_6_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 7)
    void'(lh_reg_model.Lane_7_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 8)
    void'(lh_reg_model.Lane_8_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 9)
    void'(lh_reg_model.Lane_9_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 10)
    void'(lh_reg_model.Lane_10_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 11)
    void'(lh_reg_model.Lane_11_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 12)
    void'(lh_reg_model.Lane_12_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 13)
    void'(lh_reg_model.Lane_13_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 14)
    void'(lh_reg_model.Lane_14_Status_0_CSR.Lane_Number.predict(lane_num));
  else if (lane_num == 15)
    void'(lh_reg_model.Lane_15_Status_0_CSR.Lane_Number.predict(lane_num));

endtask : update_ls0_lane_num_field



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_ls0_8b_10b_dec_err_field
/// Description : This method updates the 8B/10B decoding errors field in the LaneN_Status_0 CSR,
/// based on the invalid_cg_cnt.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_ls0_8b_10b_dec_err_field();

  forever begin //{

    @(invalid_cg_cnt);

    if (invalid_cg_cnt == 0)
      continue;

    if (lane_num == 0)
      void'(lh_reg_model.Lane_0_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 1)
      void'(lh_reg_model.Lane_1_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 2)
      void'(lh_reg_model.Lane_2_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 3)
      void'(lh_reg_model.Lane_3_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 4)
      void'(lh_reg_model.Lane_4_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 5)
      void'(lh_reg_model.Lane_5_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 6)
      void'(lh_reg_model.Lane_6_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 7)
      void'(lh_reg_model.Lane_7_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 8)
      void'(lh_reg_model.Lane_8_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 9)
      void'(lh_reg_model.Lane_9_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 10)
      void'(lh_reg_model.Lane_10_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 11)
      void'(lh_reg_model.Lane_11_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 12)
      void'(lh_reg_model.Lane_12_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 13)
      void'(lh_reg_model.Lane_13_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 14)
      void'(lh_reg_model.Lane_14_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));
    else if (lane_num == 15)
      void'(lh_reg_model.Lane_15_Status_0_CSR.lane_8B_10B_decoding_errors.predict(invalid_cg_cnt));

  end //}

endtask : update_ls0_8b_10b_dec_err_field



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_ls0_rcvr_pol_field
/// Description : This method updates the receiver input inverted field in the LaneN_Status_0 CSR,
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_ls0_rcvr_pol_field();

  ls0_rcvr_pol_field_updated = 1;

  if (lane_num == 0)
    void'(lh_reg_model.Lane_0_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 1)
    void'(lh_reg_model.Lane_1_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 2)
    void'(lh_reg_model.Lane_2_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 3)
    void'(lh_reg_model.Lane_3_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 4)
    void'(lh_reg_model.Lane_4_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 5)
    void'(lh_reg_model.Lane_5_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 6)
    void'(lh_reg_model.Lane_6_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 7)
    void'(lh_reg_model.Lane_7_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 8)
    void'(lh_reg_model.Lane_8_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 9)
    void'(lh_reg_model.Lane_9_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 10)
    void'(lh_reg_model.Lane_10_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 11)
    void'(lh_reg_model.Lane_11_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 12)
    void'(lh_reg_model.Lane_12_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 13)
    void'(lh_reg_model.Lane_13_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 14)
    void'(lh_reg_model.Lane_14_Status_0_CSR.Receiver_input_inverted.predict(1));
  else if (lane_num == 15)
    void'(lh_reg_model.Lane_15_Status_0_CSR.Receiver_input_inverted.predict(1));

endtask : update_ls0_rcvr_pol_field



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_other_ls0_fields
/// Description : This method updates the remaining fields in the LaneN_Status_0 CSR, such as
/// lane_ready, lane_sync and receiver_trained.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_other_ls0_fields();

  if (lane_num == 0)
  begin //{
    void'(lh_reg_model.Lane_0_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_0_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_0_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 1)
  begin //{
    void'(lh_reg_model.Lane_1_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_1_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_1_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 2)
  begin //{
    void'(lh_reg_model.Lane_2_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_2_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_2_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 3)
  begin //{
    void'(lh_reg_model.Lane_3_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_3_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_3_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 4)
  begin //{
    void'(lh_reg_model.Lane_4_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_4_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_4_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 5)
  begin //{
    void'(lh_reg_model.Lane_5_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_5_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_5_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 6)
  begin //{
    void'(lh_reg_model.Lane_6_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_6_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_6_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 7)
  begin //{
    void'(lh_reg_model.Lane_7_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_7_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_7_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 8)
  begin //{
    void'(lh_reg_model.Lane_8_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_8_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_8_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 9)
  begin //{
    void'(lh_reg_model.Lane_9_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_9_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_9_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 10)
  begin //{
    void'(lh_reg_model.Lane_10_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_10_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_10_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 11)
  begin //{
    void'(lh_reg_model.Lane_11_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_11_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_11_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 12)
  begin //{
    void'(lh_reg_model.Lane_12_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_12_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_12_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 13)
  begin //{
    void'(lh_reg_model.Lane_13_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_13_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_13_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 14)
  begin //{
    void'(lh_reg_model.Lane_14_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_14_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_14_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}
  else if (lane_num == 15)
  begin //{
    void'(lh_reg_model.Lane_15_Status_0_CSR.Receiver_lane_ready.predict(lh_trans.lane_ready[lane_num]));
    void'(lh_reg_model.Lane_15_Status_0_CSR.Receiver_lane_sync.predict(lh_trans.lane_sync[lane_num]));
    void'(lh_reg_model.Lane_15_Status_0_CSR.Receiver_trained.predict(lh_trans.rcvr_trained[lane_num]));
  end //}

endtask : update_other_ls0_fields



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_ls1_reg
/// Description : This method updates the LaneN_Status_1 CSR.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_ls1_reg();

  if (lane_num == 0)
    void'(lh_reg_model.Lane_0_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 1)
    void'(lh_reg_model.Lane_1_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 2)
    void'(lh_reg_model.Lane_2_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 3)
    void'(lh_reg_model.Lane_3_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 4)
    void'(lh_reg_model.Lane_4_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 5)
    void'(lh_reg_model.Lane_5_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 6)
    void'(lh_reg_model.Lane_6_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 7)
    void'(lh_reg_model.Lane_7_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 8)
    void'(lh_reg_model.Lane_8_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 9)
    void'(lh_reg_model.Lane_9_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 10)
    void'(lh_reg_model.Lane_10_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 11)
    void'(lh_reg_model.Lane_11_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 12)
    void'(lh_reg_model.Lane_12_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 13)
    void'(lh_reg_model.Lane_13_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 14)
    void'(lh_reg_model.Lane_14_Status_1_CSR.predict(lane_status_1_reg_val));
  else if (lane_num == 15)
    void'(lh_reg_model.Lane_15_Status_1_CSR.predict(lane_status_1_reg_val));

endtask : update_ls1_reg



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : sixty_sevenb_sixty_fourb_decode
/// Description : Decode method for GEN3.0. It decodes the received 67bit data into 64bit data.
/// If 'type' field is '1', then it is decoded as DATA codeword, else it is decoded as CONTROL
/// codeword. If the received codeword is a control codeword, then based on the 'cc_type' and the 
/// following 4 bits, it is decoded to identify the control codeword type, whether it is SKIP_MARKER / 
/// LANE_CHECK / SKIP / DECSR_SEED / STATUS_CNTL / CSB / CSE / CSEB. If none of the control codeword
/// decoding matches, then it is marked as invalid codeword. The decoded information is assigned to
/// the respective fields of the lane data instance which will be used by the higher level components.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::sixty_sevenb_sixty_fourb_decode();

  if (lane_data_ins.brc3_cg[2])
  begin //{ 
    lane_data_ins.brc3_type = 1; // Data codeword
    lane_data_ins.brc3_cntl_cw_type = DATA;
  end //}
  else
  begin //{

    lane_data_ins.brc3_type = 0; // Control codeword

    lane_data_ins.brc3_cc_type = lane_data_ins.brc3_cg[33:34];

    if (lane_data_ins.brc3_cc_type == 2'b00 && lane_data_ins.brc3_cg[35:38] == 4'b1011)
      lane_data_ins.brc3_cntl_cw_type = SKIP_MARKER;
    else if (lane_data_ins.brc3_cc_type == 2'b00 && lane_data_ins.brc3_cg[35:38] == 4'b1100)
      lane_data_ins.brc3_cntl_cw_type = LANE_CHECK;
    else if (lane_data_ins.brc3_cc_type == 2'b00 && lane_data_ins.brc3_cg[35:38] == 4'b1101)
      lane_data_ins.brc3_cntl_cw_type = DESCR_SEED;
    else if (lane_data_ins.brc3_cc_type == 2'b00 && lane_data_ins.brc3_cg[35:38] == 4'b1110)
      lane_data_ins.brc3_cntl_cw_type = SKIP;
    else if (lane_data_ins.brc3_cc_type == 2'b00 && lane_data_ins.brc3_cg[35:38] == 4'b1111)
      lane_data_ins.brc3_cntl_cw_type = STATUS_CNTL;
    else if (lane_data_ins.brc3_cc_type == 2'b01)
      lane_data_ins.brc3_cntl_cw_type = CSB;
    else if (lane_data_ins.brc3_cc_type == 2'b10)
      lane_data_ins.brc3_cntl_cw_type = CSE;
    else if (lane_data_ins.brc3_cc_type == 2'b11)
      lane_data_ins.brc3_cntl_cw_type = CSEB;
    else
      lane_data_ins.brc3_cntl_cw_type = INVALID_CW;

  end //}

  lane_data_ins.brc3_cw = lane_data_ins.brc3_cg[3:66];

  if (~bfm_or_mon)
  begin //{
    lc_cw_bip_calc_method(); // Temp comment. Need to uncomment once it is implemented in tx path.
  end //}
//  if (lane_data_ins.brc3_type)
//    `uvm_info("SRIO_LANE_HANDLER : GEN3 DECODE INFO", $sformatf("LANE NUM : %0d Data codeword received. Value is %0h", lane_num, lane_data_ins.brc3_cw), UVM_LOW)
//if (~bfm_or_mon && ~mon_type)
//    `uvm_info("SRIO_LANE_HANDLER : GEN3 DECODE INFO", $sformatf("LANE NUM : %0d Control codeword received. brc3_cc_type is %0h, brc3_cntl_cw_type is %0s, brc3_cw is %0h, brc3_cg is %0h", lane_num, lane_data_ins.brc3_cc_type, lane_data_ins.brc3_cntl_cw_type.name(), lane_data_ins.brc3_cw, lane_data_ins.brc3_cg), UVM_LOW)

endtask : sixty_sevenb_sixty_fourb_decode




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_data_descramble
/// Description : GEN3.0 descrambler is initialized by the receiving DESCR_SEED control codeword.
/// The first DESCR_SEED control codeword of the DESCR_SEED ordered sequence is used to initilalize
/// the descrambler lfsr, and the following DESCR_SEED codeword of the same ordered sequence is used
/// to check if the descrambler is in sync or not. Once the descrmabler is in sync, before descrambling
/// the data, the descrambler lfsr is stored in a temporary variable and it is shifted 58 times to get
/// the next lfsr value. Then, the current lfsr, and 6 bits from the shifted lfsr are used together
/// to descramble the received codeword. Finally, the current lfsr is shifted 64 times to get the new
/// lfsr seed to descramble the next data.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_data_descramble();
  bit [0:57] lcl_cpy_to_chk;				///< Holds the shifted value of GEN3.0 Descrambler LFSR

  if (lane_data_ins.brc3_cntl_cw_type == SKIP)
  begin //{

    sync_sm_descr_sync = 0;
    sync_sm_descr_err = 0;

    return;

  end //}

  if (lane_data_ins.brc3_cntl_cw_type == DESCR_SEED && descr_seed_cntl_cw_cnt == 0)
  begin //{

    lcl_cpy_to_chk=gen3_descr_lfsr;
    gen3_descr_lfsr = {lane_data_ins.brc3_cw[0:29], lane_data_ins.brc3_cw[36:63]};
    descr_seed_cntl_cw_cnt++;
     if(gen3_descr_lfsr!=lcl_cpy_to_chk && lh_trans.port_initialized)
      `uvm_error("SRIO_PL_LANE_HANDLER : GEN3_DESCRAMBLER", $sformatf(" Spec reference 5.5.4. Descrambler lfsr does not match received seed.Expected:%x Actual:%x",lcl_cpy_to_chk,gen3_descr_lfsr))

    sync_sm_descr_sync = 0;
    sync_sm_descr_err = 0;

  end //}
  else if (lane_data_ins.brc3_cntl_cw_type == DESCR_SEED && descr_seed_cntl_cw_cnt == 1)
  begin //{

    temp_gen3_descr_lfsr = {lane_data_ins.brc3_cw[0:29], lane_data_ins.brc3_cw[36:63]};

    if (temp_gen3_descr_lfsr == gen3_descr_lfsr)
    begin //{
      descr_in_sync = 1;
      sync_sm_descr_sync = 1;
      sync_sm_descr_err = 0;
    end //}
    else
    begin //{

      sync_sm_descr_sync = 0;
      sync_sm_descr_err = 1;

      if (~lh_trans.ies_state && lh_trans.link_initialized && descr_in_sync)
      begin //{
        lh_trans.ies_state = 1;
        lh_trans.ies_cause_value = 7;
        //$display($time, " 10. Vaidhy : gen3 ies_state set here");
      end //}

      descr_in_sync = 0;

      if (~bfm_or_mon)
      begin //{
        update_error_detect_csr("DESCR_SYNC_LOSS");
      end //}

    end //}

    descr_seed_cntl_cw_cnt = 0;

  end //}
  else if (lane_data_ins.brc3_cntl_cw_type != DESCR_SEED && descr_seed_cntl_cw_cnt == 1)
  begin //{

    sync_sm_descr_sync = 0;
    sync_sm_descr_err = 1;

    if (~lh_trans.ies_state && lh_trans.link_initialized && descr_in_sync)
    begin //{
      lh_trans.ies_state = 1;
      lh_trans.ies_cause_value = 7;
      //$display($time, " 11. Vaidhy : gen3 ies_state set here");
    end //}

    descr_in_sync = 0;
    
    descr_seed_cntl_cw_cnt = 0;

    if (~bfm_or_mon)
    begin //{
      update_error_detect_csr("DESCR_SYNC_LOSS");
    end //}

  end //}
  else if (lane_data_ins.brc3_cntl_cw_type != DESCR_SEED && descr_seed_cntl_cw_cnt == 0)
  begin //{

    sync_sm_descr_sync = 0;
    sync_sm_descr_err = 0;

    if (descr_in_sync)
    begin //{

      if (lane_data_ins.brc3_type || (~lane_data_ins.brc3_type && lane_data_ins.brc3_cc_type != 2'b00))
      begin //{

        temp_gen3_descr_lfsr = gen3_descr_lfsr;

        shift_gen3_descr_lfsr(58, temp_gen3_descr_lfsr);
	temp_gen3_descr_lfsr = gen3_shifted_lfsr;

	for (int bit_rev=0; bit_rev<58; bit_rev++)
	begin //{
	  reversed_gen3_descr_lfsr[bit_rev] = gen3_descr_lfsr[bit_rev];
	  reversed_temp_gen3_descr_lfsr[bit_rev] = temp_gen3_descr_lfsr[bit_rev];
	end //}

        lane_data_ins.brc3_cw = {reversed_gen3_descr_lfsr, reversed_temp_gen3_descr_lfsr[57:52]} ^ lane_data_ins.brc3_cw; // data descrambling logic.

        if(~lane_data_ins.brc3_type && lane_data_ins.brc3_cc_type != 2'b00)
         lane_data_ins.brc3_cw[30:31]=lane_data_ins.brc3_cc_type ;
      end //}

    end //}

  end //}

  shift_gen3_descr_lfsr(64, gen3_descr_lfsr);
  gen3_descr_lfsr = gen3_shifted_lfsr;

  //if (~bfm_or_mon && ~mon_type && lane_num <= 1)
  //  `uvm_info("SRIO_LANE_HANDLER : GEN3 DESCR INFO", $sformatf("LANE NUM : %0d brc3_cw is %0h", lane_num, lane_data_ins.brc3_cw), UVM_LOW)

endtask : gen3_data_descramble




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : shift_gen3_descr_lfsr
/// Description : This method is called by the gen3_data_descramble method. As per the gen3_data_descramble
/// logic, the current lfsr is shifted 58 times through a temporary lfsr variable, and finally at the
/// end of descramble logic, the current lfsr is shifted 64 times to get the new lfsr seed value. To
/// control this lfsr shift count, the integer variable shift_count is used in the method's argument.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::shift_gen3_descr_lfsr(int shift_count, bit [0:57] gen3_lfsr);

  bit lfsr_out_bit;
  bit lfsr_bit39;
  bit [0:57] lfsr_bit0_56;
  bit [0:57] local_temp_gen3_lfsr;
  int iter;

  local_temp_gen3_lfsr = gen3_lfsr;

  repeat(shift_count) begin //{

    lfsr_out_bit = local_temp_gen3_lfsr[57];
    lfsr_bit39 = local_temp_gen3_lfsr[38];
    lfsr_bit0_56 = local_temp_gen3_lfsr;
    local_temp_gen3_lfsr = {lfsr_out_bit ^ lfsr_bit39, lfsr_bit0_56[0:56]};

  end //}

  gen3_shifted_lfsr = local_temp_gen3_lfsr;

endtask : shift_gen3_descr_lfsr




//////////////////////////////////////////////////////////////////////////////////////////
/// Name : status_cntl_os_check_method
/// Description : This method checks the completeness of STATUS/CONTROL ordered sequence.
/// It also triggers the gen3_cw_training_method.
//////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::status_cntl_os_check_method();

  int rv;

  // It is enough to check the CW training logic in the first STATUS_CNTL CW of the
  // STATUS_CONTROL Ordered sequence. Thus, using the lh_status_cntl_cw_cnt to ignore
  // the CW training check in the 2nd STATUS_CNTL CW of the ordered sequence. Any
  // errors in the received ordered sequence will be taken care in the rx data handler
  // block when the corresponding ordered sequence check is performed.
  if (lane_data_ins.brc3_cntl_cw_type == STATUS_CNTL && lh_status_cntl_cw_cnt == 0 && lh_trans.lane_sync[lane_num])
  begin //{
  
    if (~lh_trans.lane_trained[lane_num])
      gen3_cw_training_method();

    lh_status_cntl_cw_cnt++;
    prev_status_cntl_cw = lane_data_ins.brc3_cw;

    if (~bfm_or_mon)
    begin //{

      rv = 29;
      for (int cwb=0; cwb<30; cwb++)
      begin //{
        ls2_reg_val[rv] = lane_data_ins.brc3_cw[cwb];
	rv--;
      end //}

      rv = 19;
      for (int cwb=36; cwb<56; cwb++)
      begin //{
        ls3_reg_val[rv] = lane_data_ins.brc3_cw[cwb];
	rv--;
      end //}

      update_ls2_reg();
      update_ls3_reg();

    end //}
  
  end //}
  else if (lane_data_ins.brc3_cntl_cw_type == STATUS_CNTL && lh_status_cntl_cw_cnt == 1)
  begin //{
  
    lh_status_cntl_cw_cnt = 0;
  
    if (prev_status_cntl_cw != lane_data_ins.brc3_cw && ~bfm_or_mon)
    begin //{
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
      `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_DIFFERENT_SC_CW_IN_SC_OS_CHECK", $sformatf(" Spec reference 5.5.3.5. Status-control control codewords in the same STATUS_CNTL ordered sequence are different. First status control codeword is %0h, Second status control codeword is %0h", prev_status_cntl_cw, lane_data_ins.brc3_cw))
    end //}
    else if (~bfm_or_mon) // if proper sc os is received.
    begin //{
      if (lane_data_ins.brc3_cw[54] || lane_data_ins.brc3_cw[55])
      begin //{
        lh_common_mon_trans.sc_os_cnt[mon_type]++;
      end //}
    end //}
  
  end //}
  else if (lane_data_ins.brc3_cntl_cw_type != STATUS_CNTL && lh_status_cntl_cw_cnt == 1 && ~bfm_or_mon)
  begin //{

    if (~lh_trans.ies_state && lh_trans.link_initialized)
    begin //{
      lh_trans.ies_state = 1;
      lh_trans.ies_cause_value = 31;
    //$display($time, " 10. Vaidhy : ies_state set here");
    end //}
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
    `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_INCOMPLETE_SC_OS_CHECK", $sformatf(" Spec reference 5.8.2. Incomplete STATUS_CNTL ordered sequence detected in IDLE3. brc3_cw_type is %0s", lane_data_ins.brc3_cntl_cw_type.name()))

    lh_status_cntl_cw_cnt = 0;
  
  end //}

endtask : status_cntl_os_check_method




/////////////////////////////////////////////////////////////////////////////////
/// Name : descr_seed_os_check_method
/// Description : This method checks the completeness of SEED ordered sequence.
/////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::descr_seed_os_check_method();

  if (lane_data_ins.brc3_cntl_cw_type == DESCR_SEED && lh_descr_seed_cw_cnt == 0 && lh_trans.lane_sync[lane_num])
  begin //{

    lh_descr_seed_cw_cnt++;
  
  end //}
  else if (lh_descr_seed_cw_cnt == 1 && lane_data_ins.brc3_cntl_cw_type != DESCR_SEED && ~bfm_or_mon)
  begin //{

    if (~lh_trans.ies_state && lh_trans.link_initialized)
    begin //{
      lh_trans.ies_state = 1;
      lh_trans.ies_cause_value = 31;
    //$display($time, " 10. Vaidhy : ies_state set here");
    end //}
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
    `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_INCOMPLETE_DS_OS_CHECK", $sformatf(" Spec reference 5.8.1. Incomplete DESCR_SEED ordered sequence detected in IDLE3. brc3_cw_type is %0s", lane_data_ins.brc3_cntl_cw_type.name()))

    lh_descr_seed_cw_cnt = 0;

  end //}
  else if (lh_descr_seed_cw_cnt == 1 && lane_data_ins.brc3_cntl_cw_type == DESCR_SEED)
  begin //{

    lh_descr_seed_cw_cnt = 0;

  end //}

endtask : descr_seed_os_check_method





/////////////////////////////////////////////////////////////////////////////////
/// Name : skip_os_check_method
/// Description : This method checks the completeness of SKIP ordered sequence.
/////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::skip_os_check_method();

  if (lane_data_ins.brc3_cntl_cw_type == SKIP_MARKER && lh_skip_os_cw_cnt == 0 && lh_trans.lane_sync[lane_num])
  begin //{

    skip_marker_cw_fixed_value_check();
    lh_skip_os_cw_cnt++;
  
  end //}
  else if (lh_skip_os_cw_cnt == 0 && lane_data_ins.brc3_cntl_cw_type == SKIP && ~bfm_or_mon)
  begin //{

    if (~lh_trans.ies_state && lh_trans.link_initialized)
    begin //{
      lh_trans.ies_state = 1;
      lh_trans.ies_cause_value = 31;
    //$display($time, " 10. Vaidhy : ies_state set here");
    end //}
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
    `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_SKIP_CW_IN_NON_SKIP_OS_CHECK", $sformatf(" Spec reference 5.8.3. SKIP control codeword received in other than skip ordered sequence"))

  end //}
  else if (lh_skip_os_cw_cnt == 0 && lane_data_ins.brc3_cntl_cw_type == LANE_CHECK && ~bfm_or_mon)
  begin //{

    if (~lh_trans.ies_state && lh_trans.link_initialized)
    begin //{
      lh_trans.ies_state = 1;
      lh_trans.ies_cause_value = 31;
    //$display($time, " 10. Vaidhy : ies_state set here");
    end //}
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
    `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_LC_CW_IN_NON_SKIP_OS_CHECK", $sformatf(" Spec reference 5.8.3. LANE_CHECK control codeword received in other than skip ordered sequence"))

  end //}
  else if (lh_skip_os_cw_cnt == 1 && lane_data_ins.brc3_cntl_cw_type != SKIP && ~bfm_or_mon)
  begin //{

    if (~lh_trans.ies_state && lh_trans.link_initialized)
    begin //{
      lh_trans.ies_state = 1;
      lh_trans.ies_cause_value = 31;
    //$display($time, " 10. Vaidhy : ies_state set here");
    end //}
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
    `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_SKIP_CW_AFTER_SKIP_MARKER_CW_CHECK", $sformatf(" Spec reference 5.8.3. One or more SKIP control codeword has to follow SKIP_MARKER control codeword in SKIP ordered sequence of IDLE3. brc3_cw_type is %0s", lane_data_ins.brc3_cntl_cw_type.name()))

  end //}
  else if ((lh_skip_os_cw_cnt == 2 || lh_skip_os_cw_cnt == 3) && (lane_data_ins.brc3_cntl_cw_type != SKIP && lane_data_ins.brc3_cntl_cw_type != LANE_CHECK))
  begin //{
    if (~lh_trans.ies_state && lh_trans.link_initialized)
    begin //{
      lh_trans.ies_state = 1;
      lh_trans.ies_cause_value = 31;
    //$display($time, " 10. Vaidhy : ies_state set here");
    end //}

    if (~bfm_or_mon)
    begin //{
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
      `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_LC_CW_AFTER_SKIP_CW_CHECK", $sformatf(" Spec reference 5.8.3. LANE_CHECK control codeword has to follow after one or more SKIP control codewords in SKIP ordered sequence of IDLE3. brc3_cw_type is %0s", lane_data_ins.brc3_cntl_cw_type.name()))
    end //}

  end //}
  else if (lh_skip_os_cw_cnt <= 3 && lane_data_ins.brc3_cntl_cw_type == LANE_CHECK)
  begin //{

    // If LANE_CHECK control codeword is received before 3 SKIP control
    // codewords, then lh_skip_os_cw_cnt is made as 4, and assumed
    // that 3 SKIP characters had been received.
    lh_skip_os_cw_cnt = 4;

  end //}
  else if ((lh_skip_os_cw_cnt == 1 || lh_skip_os_cw_cnt == 2 || lh_skip_os_cw_cnt == 3) && lane_data_ins.brc3_cntl_cw_type == SKIP)
  begin //{
    skip_cw_fixed_value_check();
  end //}
  else if (lh_skip_os_cw_cnt == 4 && lane_data_ins.brc3_cntl_cw_type != LANE_CHECK && ~bfm_or_mon)
  begin //{

    if (~lh_trans.ies_state && lh_trans.link_initialized)
    begin //{
      lh_trans.ies_state = 1;
      lh_trans.ies_cause_value = 31;
    //$display($time, " 10. Vaidhy : ies_state set here");
    end //}
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
    `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_LC_CW_AFTER_3_SKIP_CW_CHECK", $sformatf(" Spec reference 5.8.3. LANE_CHECK control codeword has to follow after 3 SKIP control codewords in SKIP ordered sequence of IDLE3. brc3_cw_type is %0s", lane_data_ins.brc3_cntl_cw_type.name()))

  end //}
  else if ((lh_skip_os_cw_cnt == 5 || lh_skip_os_cw_cnt == 6) && (lane_data_ins.brc3_cntl_cw_type != DESCR_SEED && ~bfm_or_mon))
  begin //{

    if (~lh_trans.ies_state && lh_trans.link_initialized)
    begin //{
      lh_trans.ies_state = 1;
      lh_trans.ies_cause_value = 31;
    //$display($time, " 10. Vaidhy : ies_state set here");
    end //}
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
    `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_DS_OS_AFTER_LC_CW_CHECK", $sformatf(" Spec reference 5.8.3. DESCR_SEED ordered sequence has to follow LANE_CHECK control codeword in SKIP ordered sequence of IDLE3. brc3_cw_type is %0s", lane_data_ins.brc3_cntl_cw_type.name()))

  end //}

  if (lh_skip_os_cw_cnt == 6)
  begin //{
    lh_skip_os_cw_cnt = 0;
  end //}
  else if (lh_skip_os_cw_cnt > 0 && lane_data_ins.brc3_cntl_cw_type != SKIP_MARKER)
  begin //{
    lh_skip_os_cw_cnt++;
  end //}

endtask : skip_os_check_method




//////////////////////////////////////////////////////////////////////////////////////////////
/// Name : skip_marker_cw_fixed_value_check
/// Description : This method checks the Fixed value received in SKIP_MARKER control codeword.
//////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::skip_marker_cw_fixed_value_check();

  if (lane_data_ins.brc3_cw[0:29] != 30'h394D_E8D1 && ~bfm_or_mon)
  begin //{
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
    `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_SKIP_MARKER_FIXED_VALUE_1_CHECK", $sformatf(" Spec reference 5.5.3.1. First part of fixed value in SKIP_MARKER control codeword is different. Fixed value received is %0h. Expected  is 30'h394D_E8D1", lane_data_ins.brc3_cw[0:29]))
  end //}

  if (lane_data_ins.brc3_cw[36:63] != 28'h85E_2FA0 && ~bfm_or_mon)
  begin //{
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
    `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_SKIP_MARKER_FIXED_VALUE_2_CHECK", $sformatf(" Spec reference 5.5.3.1. Second part of fixed value in SKIP_MARKER control codeword is different. Fixed value received is %0h. Expected  is 28'h85E_2FA0", lane_data_ins.brc3_cw[36:63]))
  end //}

endtask : skip_marker_cw_fixed_value_check




///////////////////////////////////////////////////////////////////////////////////////
/// Name : skip_cw_fixed_value_check
/// Description : This method checks the Fixed value received in SKIP control codeword.
///////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::skip_cw_fixed_value_check();

  if (lane_data_ins.brc3_cw[0:29] != 30'h2E17_8BE8 && ~bfm_or_mon)
  begin //{
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
    `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_SKIP_CW_FIXED_VALUE_1_CHECK", $sformatf(" Spec reference 5.5.3.1. First part of fixed value in SKIP control codeword is different. Fixed value received is %0h. Expected  is 30'h2E17_8BE8", lane_data_ins.brc3_cw[0:29]))
  end //}

  if (lane_data_ins.brc3_cw[36:63] != 28'h537_A344 && ~bfm_or_mon)
  begin //{
      //update_error_detect_csr("INVALID_OS"); // Temp comment till the field is added in the register model.
    `uvm_error("SRIO_PL_LANE_HANDLER : IDLE3_SEQUENCE_SKIP_CW_FIXED_VALUE_2_CHECK", $sformatf(" Spec reference 5.5.3.1. Second part of fixed value in SKIP control codeword is different. Fixed value received is %0h. Expected  is 28'h537_A344", lane_data_ins.brc3_cw[36:63]))
  end //}

endtask : skip_cw_fixed_value_check




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_cw_training_method
/// Description : This method is called by the GEN3.0 logic of ser2par method.
/// Once a STATUS_CNTL codeword is received after lane_sync is achieved, this method is called to
/// decode the traning command, tap and status fields. The decoded fields are assigned to corresponding
/// variables available in the common component transaction, inorder to pass the information to the
/// transmit path of the BFM, to act accordingly based on the received training information.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_cw_training_method();

  gen3_train_data_ins = new();

  gen3_train_data_ins.xmit_equalizer_tap    = lane_data_ins.brc3_cw[41:44];
  gen3_train_data_ins.xmit_equalizer_cmd    = lane_data_ins.brc3_cw[45:47];
  gen3_train_data_ins.xmit_equalizer_status = lane_data_ins.brc3_cw[48:50];

  lh_trans.gen3_training_equalizer_tap[lane_num]    = gen3_train_data_ins.xmit_equalizer_tap;
  lh_trans.gen3_training_equalizer_cmd[lane_num]    = gen3_train_data_ins.xmit_equalizer_cmd;
  lh_trans.gen3_training_equalizer_status[lane_num] = gen3_train_data_ins.xmit_equalizer_status;

  if (gen3_train_data_ins.xmit_equalizer_cmd != 3'b000)
  begin //{
    lh_trans.gen3_training_cmd_set[lane_num] = 1;
  end //}
  else
  begin //{
    lh_trans.gen3_training_cmd_set[lane_num] = 0;
  end //}

  if (~bfm_or_mon)
  begin //{

    gen3_training_checks();

  end //}

endtask : gen3_cw_training_method



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_training_checks
/// Description : This method performs the training related checks for GEN3.0 similar to the IDLE2
/// AET checks. This method performs checks for both CW training and DME training based on the
/// training method.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_training_checks();

  if (~lh_common_mon_trans.gen3_training_cmd_outstanding[mon_type][lane_num])
  begin //{

    if (gen3_train_data_ins.xmit_equalizer_cmd != 3'b000 || ((gen3_train_data_ins.xmit_equalizer_cp1_cmd != 2'b00 || gen3_train_data_ins.xmit_equalizer_cn1_cmd != 2'b00) && lh_trans.frame_lock[lane_num]))
    begin //{

      if (lh_common_mon_trans.gen3_training_status_received[~mon_type][lane_num])
      begin //{

    	`uvm_error("SRIO_PL_LANE_HANDLER: GEN3_TRAINING_CMD_ASSERTION_CHECK", $sformatf(" Spec reference 5.10.2.2. Lane number is %0d. Transmit equalizer command shall not be assered when status is other than not_updated", lane_num))

      end //}

      if (lh_trans.frame_lock[lane_num])
      begin //{

	lh_common_mon_trans.gen3_c0_training_cmd[mon_type][lane_num] = gen3_train_data_ins.xmit_equalizer_cmd;
	lh_common_mon_trans.gen3_cp1_training_cmd[mon_type][lane_num] = gen3_train_data_ins.xmit_equalizer_cp1_cmd;
	lh_common_mon_trans.gen3_cn1_training_cmd[mon_type][lane_num] = gen3_train_data_ins.xmit_equalizer_cn1_cmd;

      end //}

      bkp_gen3_train_data_ins = new gen3_train_data_ins;
      lh_common_mon_trans.gen3_training_cmd_outstanding[mon_type][lane_num] = 1;

      if (lh_trans.lane_sync[lane_num])
        -> start_100us_cmd_timer;

    end //}

  end //}
  else
  begin //{

    if (~lh_common_mon_trans.gen3_training_status_received[~mon_type][lane_num])
    begin //{

      if (((lh_common_mon_trans.gen3_cmd_deassertion_timer_started[mon_type][lane_num] || gen3_cmd_deassertion_timer_done) && gen3_train_data_ins.xmit_equalizer_cmd == 3'b000 && lh_trans.lane_sync[lane_num]) || (lh_trans.frame_lock[lane_num] && gen3_train_data_ins.xmit_equalizer_cmd == 3'b000 && gen3_train_data_ins.xmit_equalizer_cp1_cmd == 2'b00 && gen3_train_data_ins.xmit_equalizer_cn1_cmd == 2'b00))
      begin //{

	bkp_gen3_train_data_ins = gen3_train_data_ins;
        lh_common_mon_trans.gen3_training_cmd_outstanding[mon_type][lane_num] = 0;

      end //}

      if (bkp_gen3_train_data_ins.xmit_equalizer_cmd != gen3_train_data_ins.xmit_equalizer_cmd || ((bkp_gen3_train_data_ins.xmit_equalizer_cp1_cmd != gen3_train_data_ins.xmit_equalizer_cp1_cmd || bkp_gen3_train_data_ins.xmit_equalizer_cn1_cmd != gen3_train_data_ins.xmit_equalizer_cn1_cmd) && lh_trans.frame_lock[lane_num]))
      begin //{

    	if (gen3_cmd_deassertion_timer_done && lh_trans.lane_sync[lane_num])
    	begin //{

    	  `uvm_error("SRIO_PL_LANE_HANDLER: GEN3_TRAINING_CMD_DEASSERTION_AFTER_STATUS_TIMEOUT_CHECK", $sformatf(" Spec reference 5.10.2.2. Lane number is %0d. Transmit equalizer command should be deasserted within 5us after 100us status timeout", lane_num))

    	end //}
    	else if ((~gen3_cmd_deassertion_timer_done && lh_trans.lane_sync[lane_num]) || lh_trans.frame_lock[lane_num])
    	begin //{

      	  `uvm_error("SRIO_PL_LANE_HANDLER: GEN3_TRAINING_CMD_CHANGE_BEFORE_STATUS_CHECK", $sformatf(" Spec reference 5.10.2.2. Lane number is %0d. Transmit equalizer command field shall not change before transmit equalizer status is received", lane_num))

    	end //}

      end //}

      if (bkp_gen3_train_data_ins.xmit_equalizer_tap != gen3_train_data_ins.xmit_equalizer_tap)
      begin //{

      	`uvm_error("SRIO_PL_LANE_HANDLER: GEN3_TRAINING_TAP_CHANGE_BEFORE_STATUS_CHECK", $sformatf(" Spec reference 5.10.2.2. Lane number is %0d. Transmit equalizer tap field shall not change before transmit equalizer status is received", lane_num))

      end //}

      if (gen3_cmd_deassertion_timer_done && (bkp_gen3_train_data_ins.xmit_equalizer_cmd != 0) && lh_trans.lane_sync[lane_num])
      begin //{
	// cmd deassertion timer checked only for CW training. Hence lane_sync condition added in 'if' conditions.
	// DME training doesn't specify any timers for cmd deassertion.
	bkp_gen3_train_data_ins.xmit_equalizer_cmd = 0;
      end //}

    end //}
    else
    begin //{

      if (gen3_train_data_ins.xmit_equalizer_cmd == 3'b000 && lh_trans.lane_sync[lane_num] || (gen3_train_data_ins.xmit_equalizer_cmd == 3'b000 && gen3_train_data_ins.xmit_equalizer_cp1_cmd == 2'b00 && gen3_train_data_ins.xmit_equalizer_cn1_cmd == 2'b00 && lh_trans.frame_lock[lane_num]))
      begin //{

	bkp_gen3_train_data_ins = gen3_train_data_ins;
        lh_common_mon_trans.gen3_training_cmd_outstanding[mon_type][lane_num] = 0;

      end //}
      else
      begin //{

    	if (gen3_cmd_deassertion_timer_done && lh_trans.lane_sync[lane_num])
    	begin //{

    	  `uvm_error("SRIO_PL_LANE_HANDLER: GEN3_TRAINING_CMD_DEASSERTION_AFTER_STATUS_CHECK", $sformatf(" Spec reference 5.10.2.2. Lane number is %0d. Transmit equalizer command should be deasserted within 5us of receiving status", lane_num))

    	end //}

      end //}	

    end //}

  end //}

  if (lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
  begin //{

    if ((gen3_train_data_ins.xmit_equalizer_status != 3'b000 && lh_trans.lane_sync[lane_num]) || (gen3_train_data_ins.xmit_equalizer_status != 3'b000 && gen3_train_data_ins.xmit_equalizer_cp1_status != 2'b00 && gen3_train_data_ins.xmit_equalizer_cn1_status != 2'b00 && lh_trans.frame_lock[lane_num]))
    begin //{

      lh_common_mon_trans.gen3_training_status_received[mon_type][lane_num] = 1;

      if (lh_trans.frame_lock[lane_num])
      begin //{

	if ((lh_common_mon_trans.gen3_expected_c0_training_status[mon_type][lane_num] != gen3_train_data_ins.xmit_equalizer_status) || (lh_common_mon_trans.gen3_expected_cp1_training_status[mon_type][lane_num] != gen3_train_data_ins.xmit_equalizer_cp1_status) || (lh_common_mon_trans.gen3_expected_cn1_training_status[mon_type][lane_num] != gen3_train_data_ins.xmit_equalizer_cn1_status))
	begin //{

    	  `uvm_error("SRIO_PL_LANE_HANDLER: GEN3_TRAINING_COEFF_STATUS_MISMATCH_CHECK", $sformatf(" Spec reference 802.3-2008, 72.6.10.2.4. Lane number is %0d. Expected and actual coefficient status doesn't match. Expected c0 status is %0b, Actual c0 status is %0b, Expected cp1 status is %0b, Actual cp1 status is %0b, Expected cn1 status is %0b, Actual cn1 status is %0b, ", lane_num, lh_common_mon_trans.gen3_expected_c0_training_status[mon_type][lane_num], gen3_train_data_ins.xmit_equalizer_status, lh_common_mon_trans.gen3_expected_cp1_training_status[mon_type][lane_num], gen3_train_data_ins.xmit_equalizer_cp1_status, lh_common_mon_trans.gen3_expected_cn1_training_status[mon_type][lane_num], gen3_train_data_ins.xmit_equalizer_cn1_status))

	end //}

      end //}

    end //}

  end //}
  else if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num] && lh_common_mon_trans.gen3_training_status_received[mon_type][lane_num])
  begin //{

    if ((gen3_train_data_ins.xmit_equalizer_status == 3'b000 && lh_trans.lane_sync[lane_num]) || (gen3_train_data_ins.xmit_equalizer_status == 3'b000 && gen3_train_data_ins.xmit_equalizer_cp1_status == 2'b00 && gen3_train_data_ins.xmit_equalizer_cn1_status == 2'b00 && lh_trans.frame_lock[lane_num]))
    begin //{

      lh_common_mon_trans.gen3_training_status_received[mon_type][lane_num] = 0;

    end //}

  end //}
  else if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num] && ~lh_common_mon_trans.gen3_training_status_received[mon_type][lane_num])
  begin //{

    if ((gen3_train_data_ins.xmit_equalizer_status != 3'b000 && lh_trans.lane_sync[lane_num]) || (gen3_train_data_ins.xmit_equalizer_status != 3'b000 && gen3_train_data_ins.xmit_equalizer_cp1_status != 2'b00 && gen3_train_data_ins.xmit_equalizer_cn1_status != 2'b00 && lh_trans.frame_lock[lane_num]))
    begin //{

      `uvm_error("SRIO_PL_LANE_HANDLER: GEN3_TRAINING_STATUS_WITHOUT_CMD_CHECK", $sformatf(" Spec reference 5.10.2.2. Lane number is %0d. Transmit equalizer status should not be other than not_updated when there is no active command-status handshake is outstanding", lane_num))

    end //}

  end //}

endtask : gen3_training_checks



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_cw_training_cmd_timer_method
/// Description : This method runs different timers used for GEN3.0 CW training, such as
/// ack timeout timer and command deassertion timer.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_cw_training_cmd_timer_method();

  forever
  begin //{

    wait(start_100us_cmd_timer.triggered);

    repeat(lh_config.cw_training_ack_timeout_period)
    begin //{

      if (~lh_common_mon_trans.gen3_training_status_received[~mon_type][lane_num])
        @(posedge srio_if.sim_clk);
      else
        break;

    end //}

    lh_common_mon_trans.gen3_cmd_deassertion_timer_started[mon_type][lane_num] = 1;	// 5us timer should start once the 100 us timer is completed.

    repeat(lh_config.cw_training_cmd_deassertion_period)
    begin //{

      if (lh_common_mon_trans.gen3_training_cmd_outstanding[mon_type][lane_num])
        @(posedge srio_if.sim_clk);
      else
        break;

    end //}

    lh_common_mon_trans.gen3_cmd_deassertion_timer_started[mon_type][lane_num] = 0;

    if (lh_common_mon_trans.gen3_training_cmd_outstanding[mon_type][lane_num])
    begin //{

      gen3_cmd_deassertion_timer_done = 1;

      wait (lh_common_mon_trans.gen3_training_cmd_outstanding[mon_type][lane_num] == 0);

      gen3_cmd_deassertion_timer_done = 0;

    end //}

  end //}

endtask : gen3_cw_training_cmd_timer_method



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_train_timer
/// Description : This method runs GEN3.0 training timer. Once the train_lane is set by either
/// CW training or DME trainng state machine, the gen3_training_timer is started. The timer runs till
/// it expires or till the train_lane is deasserted.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_train_timer();

  forever begin //{

    wait (lh_trans.train_lane[lane_num] == 1);

    repeat (lh_config.gen3_training_timer)
    begin //{

      if (lh_trans.train_lane[lane_num])
        @(posedge srio_if.sim_clk);
      else
        break;

    end //}

    if (lh_trans.train_lane[lane_num])
    begin //{
      lh_trans.train_timer_done[lane_num] = 1;
    end //}

  // 5 clock delay given so that train_timer_done if set, can be sampled by the
  // state machine and move the state accordingly.
    repeat(5) @(posedge srio_if.sim_clk);
    lh_trans.train_timer_done[lane_num] = 0;

    wait (lh_trans.train_lane[lane_num] == 0);

  end //}

endtask : gen3_train_timer



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_keep_alive_timer_method
/// Description : This method runs GEN3.0 keep_alive timer.
/// Once the cw training state machine enters TRAINED state, keep_alive assertion timer is started,
/// and when it expires, the keep_alive signal is asserted, which will cause the training state to
/// move to KEEP_ALIVE state. Now, the keep_alive deassertion is started, and when it expires, the
/// keep_alive signal is deasserted and the training state machine returns back to the TRAINED state.
/// At any point if the training state moves to the UNTRAINED state, then the method deasserts the
/// keep_alive signal if set and continues to wait for the TRAINED state to be reached. This method
/// runs forever.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_keep_alive_timer_method();

  forever begin //{

    wait (current_cw_train_state == TRAINED && lh_trans.current_init_state == ASYM_MODE);

    repeat (lh_config.gen3_keep_alive_assert_timer)
    begin //{

      if (~lh_trans.retrain && current_cw_train_state == TRAINED)
        @(posedge srio_if.sim_clk);
      else
        break;

    end //}

    if (~lh_trans.retrain && current_cw_train_state == TRAINED)
    begin //{
      lh_trans.keep_alive[lane_num] = 1;
    end //}

    wait (current_cw_train_state == KEEP_ALIVE || current_cw_train_state == UNTRAINED);

    if (current_cw_train_state == UNTRAINED)
    begin //{
      lh_trans.keep_alive[lane_num] = 0;
      continue;
    end //}

    repeat (lh_config.gen3_keep_alive_deassert_timer)
    begin //{

      if (~lh_trans.retrain && current_cw_train_state == KEEP_ALIVE)
        @(posedge srio_if.sim_clk);
      else
        break;

    end //}

    lh_trans.keep_alive[lane_num] = 0;

  end //}

endtask : gen3_keep_alive_timer_method



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_dme_training_commands_decode
/// Description : When a complete DME frame is received, this method decodes the control channel of
/// the frame and assigns the coefficient command and status fields. Similar to the other training
/// decode methods, this method also assigns the training information to corresponding variables
/// in the common component transaction, with which the transmit path can decide on its outbound
/// training frame.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_dme_training_commands_decode();

  forever begin //{

    wait (frame_offset_achieved == 1 && good_markers > 0);

    dme_coeff_update_status_field = complete_dme_frame[32:287];

    gen3_dme_decode(dme_coeff_update_status_field);
    decoded_dme_coeff_update_field = decoded_dme_data[0:15];
    decoded_dme_status_field = decoded_dme_data[16:31];

    gen3_train_data_ins = new();

    if (decoded_dme_coeff_update_field[13])  // preset command
    begin //{
      gen3_train_data_ins.xmit_equalizer_cmd = 3'b110;
    end //}
    else if (decoded_dme_coeff_update_field[12])  // preset command
    begin //{
      gen3_train_data_ins.xmit_equalizer_cmd = 3'b101;
    end //}
    else if (decoded_dme_coeff_update_field[3:2] == 2'b01)  // Increment and decrement encodings are interchanged in CW and DME training.
    begin //{
      gen3_train_data_ins.xmit_equalizer_cmd = 2'b10;	    // xmit_equalizer_cmd contains c0 coeff value for DME training.
    end //}
    else if (decoded_dme_coeff_update_field[3:2] == 2'b10)
    begin //{
      gen3_train_data_ins.xmit_equalizer_cmd = 2'b01;
    end //}
    else if (decoded_dme_coeff_update_field[3:2] == 2'b00)
    begin //{
      gen3_train_data_ins.xmit_equalizer_cmd = 2'b00;
    end //}

    if (decoded_dme_coeff_update_field[5:4] == 2'b01)  		// Increment and decrement encodings are interchanged in CW and DME training.
    begin //{
      gen3_train_data_ins.xmit_equalizer_cp1_cmd = 2'b10;       // xmit_equalizer_cmd contains c0 coeff value for DME training.
    end //}
    else if (decoded_dme_coeff_update_field[5:4] == 2'b10)
    begin //{
      gen3_train_data_ins.xmit_equalizer_cp1_cmd = 2'b01;
    end //}
    else if (decoded_dme_coeff_update_field[5:4] == 2'b00)
    begin //{
      gen3_train_data_ins.xmit_equalizer_cp1_cmd = 2'b00;
    end //}

    if (decoded_dme_coeff_update_field[1:0] == 2'b01)  		// Increment and decrement encodings are interchanged in CW and DME training.
    begin //{
      gen3_train_data_ins.xmit_equalizer_cn1_cmd = 2'b10;       // xmit_equalizer_cmd contains c0 coeff value for DME training.
    end //}
    else if (decoded_dme_coeff_update_field[1:0] == 2'b10)
    begin //{
      gen3_train_data_ins.xmit_equalizer_cn1_cmd = 2'b01;
    end //}
    else if (decoded_dme_coeff_update_field[1:0] == 2'b00)
    begin //{
      gen3_train_data_ins.xmit_equalizer_cn1_cmd = 2'b00;
    end //}

    //lh_trans.from_dme_rcvr_ready[lane_num] = decoded_dme_status_field[15]; // Temp comment. Need to uncomment when it is supported in tx path.
    gen3_train_data_ins.xmit_equalizer_cp1_status = decoded_dme_status_field[5:4];
    gen3_train_data_ins.xmit_equalizer_status = decoded_dme_status_field[3:2];
    gen3_train_data_ins.xmit_equalizer_cn1_status = decoded_dme_status_field[1:0];

    lh_trans.gen3_training_equalizer_tap[lane_num]    = gen3_train_data_ins.xmit_equalizer_tap;
    lh_trans.gen3_training_equalizer_cmd[lane_num]    = gen3_train_data_ins.xmit_equalizer_cmd;
    lh_trans.gen3_training_equalizer_status[lane_num] = gen3_train_data_ins.xmit_equalizer_status;

    lh_trans.gen3_training_equalizer_cp1_cmd[lane_num]    = gen3_train_data_ins.xmit_equalizer_cp1_cmd;
    lh_trans.gen3_training_equalizer_cn1_cmd[lane_num]    = gen3_train_data_ins.xmit_equalizer_cn1_cmd;

    lh_trans.gen3_training_equalizer_cp1_status[lane_num]    = gen3_train_data_ins.xmit_equalizer_cp1_status;
    lh_trans.gen3_training_equalizer_cn1_status[lane_num]    = gen3_train_data_ins.xmit_equalizer_cn1_status;

    if (gen3_train_data_ins.xmit_equalizer_cmd != 3'b000)
    begin //{
      lh_trans.gen3_training_cmd_set[lane_num] = 1;
    end //}
    else
    begin //{
      lh_trans.gen3_training_cmd_set[lane_num] = 0;
    end //}

    if (gen3_train_data_ins.xmit_equalizer_cp1_cmd != 2'b00)
    begin //{
      lh_trans.gen3_training_cp1_cmd_set[lane_num] = 1;
    end //}
    else
    begin //{
      lh_trans.gen3_training_cp1_cmd_set[lane_num] = 0;
    end //}

    if (gen3_train_data_ins.xmit_equalizer_cn1_cmd != 2'b00)
    begin //{
      lh_trans.gen3_training_cn1_cmd_set[lane_num] = 1;
    end //}
    else
    begin //{
      lh_trans.gen3_training_cn1_cmd_set[lane_num] = 0;
    end //}

    if (~bfm_or_mon && ~lh_trans.lane_trained[lane_num])
    begin //{

      gen3_training_checks();

    end //}

    wait (frame_offset_achieved == 0 || bad_markers > 0);

  end //}

endtask : gen3_dme_training_commands_decode



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_dme_decode
/// Description : This is the decoder method for differential manchester encoded control channel of
/// a training frame. Based on the protocol, if the 8-bit data has a mid-cell data transition, then
/// it is decoded as a '1' or else it is decoded as a '0'.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_dme_decode(bit [0:255] dme_data);

  int decoded_data_bit;
  bit [0:7] temp_dme_byte;

  decoded_data_bit = 0;

  for (int dbs=0; dbs<255; dbs=dbs+8)
  begin //{

    temp_dme_byte = dme_data[dbs+:8];

    if (temp_dme_byte[0:3] == ~temp_dme_byte[4:7])
      decoded_dme_data[decoded_data_bit] = 1;
    else if (temp_dme_byte[0:3] == temp_dme_byte[4:7])
      decoded_dme_data[decoded_data_bit] = 0;
    else
    begin //{
      `uvm_warning("SRIO_PL_LANE_HANDLER : DME_DATA_DECODE", $sformatf(" Spec reference 802.3-2008, 72.6.10.2.2. Lane number %0d : DME data not encoded properly. Transition shall happen on either cell boundary or half-cell boundary. Bit position %0d to %0d, 8 bit data received is %0h", lane_num, dbs, dbs+8, temp_dme_byte))
    end //}

    decoded_data_bit++;
    
  end //}

endtask : gen3_dme_decode



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_c0_coeff_update_sm
/// Description : This is the coefficient update state machine for main tap C0. The state machine
/// is defined in the 802.3-2008 specification.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_c0_coeff_update_sm();

#1;
  if (~srio_if.srio_rst_n)
  begin //{

    current_c0_coeff_update_state = NOT_UPDATED;
    // questasim and vcs doesn't work properly on associatuve array methods
    // Hence, a work-around is done here by setting the array values to 1 and
    // then clearing it immediately.
    lh_trans.gen3_training_cmd_set[lane_num] = 1;
    lh_trans.gen3_training_cmd_set[lane_num] = 0;

    lh_trans.gen3_training_cp1_cmd_set[lane_num] = 1;
    lh_trans.gen3_training_cp1_cmd_set[lane_num] = 0;

    lh_trans.gen3_training_cn1_cmd_set[lane_num] = 1;
    lh_trans.gen3_training_cn1_cmd_set[lane_num] = 0;

    if (~bfm_or_mon)
    begin //{

      lh_common_mon_trans.gen3_c0_training_cmd[mon_type][lane_num] = 1;
      lh_common_mon_trans.gen3_c0_training_cmd[mon_type][lane_num] = 0;

      lh_common_mon_trans.gen3_cp1_training_cmd[mon_type][lane_num] = 1;
      lh_common_mon_trans.gen3_cp1_training_cmd[mon_type][lane_num] = 0;

      lh_common_mon_trans.gen3_cn1_training_cmd[mon_type][lane_num] = 1;
      lh_common_mon_trans.gen3_cn1_training_cmd[mon_type][lane_num] = 0;

      lh_common_mon_trans.gen3_expected_c0_training_status[mon_type][lane_num] = 1;
      lh_common_mon_trans.gen3_expected_c0_training_status[mon_type][lane_num] = 0;

      lh_common_mon_trans.gen3_expected_cp1_training_status[mon_type][lane_num] = 1;
      lh_common_mon_trans.gen3_expected_cp1_training_status[mon_type][lane_num] = 0;

      lh_common_mon_trans.gen3_expected_cn1_training_status[mon_type][lane_num] = 1;
      lh_common_mon_trans.gen3_expected_cn1_training_status[mon_type][lane_num] = 0;

    end //}

    if (bfm_or_mon)
    begin //{
      c0_preset_value = lh_config.bfm_dme_training_c0_preset_value;
      c0_init_value = lh_config.bfm_dme_training_c0_init_value;
      c0_max_limit = lh_config.bfm_dme_training_c0_max_value;
      c0_min_limit = lh_config.bfm_dme_training_c0_min_value;
    end //}
    else if (mon_type && lh_env_config.srio_tx_mon_if == DUT)
    begin //{
      c0_preset_value = lh_config.bfm_dme_training_c0_preset_value;
      c0_init_value = lh_config.bfm_dme_training_c0_init_value;
      c0_max_limit = lh_config.bfm_dme_training_c0_max_value;
      c0_min_limit = lh_config.bfm_dme_training_c0_min_value;
    end //}
    else if (mon_type && lh_env_config.srio_tx_mon_if == BFM)
    begin //{
      c0_preset_value = lh_config.lp_dme_training_c0_preset_value;
      c0_init_value = lh_config.lp_dme_training_c0_init_value;
      c0_max_limit = lh_config.lp_dme_training_c0_max_value;
      c0_min_limit = lh_config.lp_dme_training_c0_min_value;
    end //}
    else if (~mon_type && lh_env_config.srio_rx_mon_if == DUT)
    begin //{
      c0_preset_value = lh_config.bfm_dme_training_c0_preset_value;
      c0_init_value = lh_config.bfm_dme_training_c0_init_value;
      c0_max_limit = lh_config.bfm_dme_training_c0_max_value;
      c0_min_limit = lh_config.bfm_dme_training_c0_min_value;
    end //}
    else if (~mon_type && lh_env_config.srio_rx_mon_if == BFM)
    begin //{
      c0_preset_value = lh_config.lp_dme_training_c0_preset_value;
      c0_init_value = lh_config.lp_dme_training_c0_init_value;
      c0_max_limit = lh_config.lp_dme_training_c0_max_value;
      c0_min_limit = lh_config.lp_dme_training_c0_min_value;
    end //}

    if (~bfm_or_mon)
      current_c0_coeff_update_state_q.push_back(current_c0_coeff_update_state);

  end //}

  forever
  begin //{

    wait (lh_trans.frame_lock[lane_num] == 1);

    @(negedge dme_frame_divide_clk or negedge srio_if.srio_rst_n);

    if (~srio_if.srio_rst_n || lh_trans.mr_restart_training)
    begin //{

      prev_c0_coeff_update_state = current_c0_coeff_update_state;

      current_c0_coeff_update_state = NOT_UPDATED;
      lh_trans.gen3_c0_coeff_status[lane_num] = 2'b00;

      if (~bfm_or_mon)
      begin //{
        lh_common_mon_trans.gen3_expected_c0_training_status[~mon_type][lane_num] = 2'b00;
      end //}

      if (~bfm_or_mon && prev_c0_coeff_update_state != current_c0_coeff_update_state)
        current_c0_coeff_update_state_q.push_back(current_c0_coeff_update_state);

    end //}
    else
    begin //{

      //`uvm_info("SRIO_LANE_HANDLER : GEN3_CW_TRAIN_SM", $sformatf(" lane_trained[%0d] is %0d Present cw train state is %0s", lane_num, lh_trans.lane_trained[lane_num], current_dme_train_state.name()), UVM_LOW)

      prev_c0_coeff_update_state = current_c0_coeff_update_state;

      case (current_c0_coeff_update_state)

	NOT_UPDATED : begin //{

      			lh_trans.gen3_c0_coeff_status[lane_num] = 2'b00;

      			if (~bfm_or_mon)
      			begin //{

      			  lh_common_mon_trans.gen3_expected_c0_training_status[mon_type][lane_num] = 2'b00;

		      	  if (lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      	  begin //{
      		      	    current_c0_coeff_update_state = UPDATE_COEFF;
		      	  end //}

      			end //}
			else
			begin //{

		      	  if (lh_trans.gen3_training_cmd_set[lane_num])
		      	  begin //{
      		      	    current_c0_coeff_update_state = UPDATE_COEFF;
		      	  end //}

			end //}

		      end //}

	UPDATE_COEFF : begin //{

      			if (~bfm_or_mon)
      			begin //{

		      	  if (lh_common_mon_trans.gen3_c0_training_cmd[~mon_type][lane_num] == 3'b110)	// preset
		      	  begin //{
      		      	    new_c0_coeff = c0_preset_value;
		      	  end //}
		      	  else if (lh_common_mon_trans.gen3_c0_training_cmd[~mon_type][lane_num] == 3'b101) // Initialize
		      	  begin //{
      		      	    new_c0_coeff = c0_init_value;
		      	  end //}
		      	  else if (lh_common_mon_trans.gen3_c0_training_cmd[~mon_type][lane_num] == 3'b010) // Increment
		      	  begin //{
      		      	    new_c0_coeff = (new_c0_coeff < c0_max_limit) ? new_c0_coeff+1 : c0_max_limit;
		      	  end //}
		      	  else if (lh_common_mon_trans.gen3_c0_training_cmd[~mon_type][lane_num] == 3'b001) // decrement
		      	  begin //{
      		      	    new_c0_coeff = (new_c0_coeff > c0_min_limit) ? new_c0_coeff-1 : c0_min_limit;
		      	  end //}

      			end //}
			else
			begin //{


		      	  if (lh_trans.gen3_training_equalizer_cmd[lane_num] == 3'b110)	// preset
		      	  begin //{
      		      	    new_c0_coeff = c0_preset_value;
		      	  end //}
		      	  else if (lh_trans.gen3_training_equalizer_cmd[lane_num] == 3'b101) // Initialize
		      	  begin //{
      		      	    new_c0_coeff = c0_init_value;
		      	  end //}
		      	  else if (lh_trans.gen3_training_equalizer_cmd[lane_num] == 3'b010) // Increment
		      	  begin //{
      		      	    new_c0_coeff = (new_c0_coeff < c0_max_limit) ? new_c0_coeff+1 : c0_max_limit;
		      	  end //}
		      	  else if (lh_trans.gen3_training_equalizer_cmd[lane_num] == 3'b001) // decrement
		      	  begin //{
      		      	    new_c0_coeff = (new_c0_coeff > c0_min_limit) ? new_c0_coeff-1 : c0_min_limit;
		      	  end //}

			end //}

			if (new_c0_coeff >= c0_max_limit)
			  current_c0_coeff_update_state = MAXIMUM;
			else if ((new_c0_coeff > c0_min_limit) && (new_c0_coeff < c0_max_limit))
			  current_c0_coeff_update_state = UPDATED;
			else if (new_c0_coeff <= c0_max_limit)
			  current_c0_coeff_update_state = MINIMUM;

		      end //}

	MAXIMUM : begin //{

      		    lh_trans.gen3_c0_coeff_status[lane_num] = 2'b11;

      		    if (~bfm_or_mon)
      		    begin //{

      		      lh_common_mon_trans.gen3_expected_c0_training_status[mon_type][lane_num] = 2'b11;

		      if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      begin //{
      		        current_c0_coeff_update_state = NOT_UPDATED;
		      end //}

      		    end //}
		    else
		    begin //{

		      if (~lh_trans.gen3_training_cmd_set[lane_num])
		      begin //{
      		        current_c0_coeff_update_state = NOT_UPDATED;
		      end //}

		    end //}

	    	  end //}

	UPDATED : begin //{

      		    lh_trans.gen3_c0_coeff_status[lane_num] = 2'b01;

      		    if (~bfm_or_mon)
      		    begin //{

      		      lh_common_mon_trans.gen3_expected_c0_training_status[mon_type][lane_num] = 2'b01;

		      if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      begin //{
      		        current_c0_coeff_update_state = NOT_UPDATED;
		      end //}

      		    end //}
		    else
		    begin //{

		      if (~lh_trans.gen3_training_cmd_set[lane_num])
		      begin //{
      		        current_c0_coeff_update_state = NOT_UPDATED;
		      end //}

		    end //}

	    	  end //}

	MINIMUM : begin //{

      		    lh_trans.gen3_c0_coeff_status[lane_num] = 2'b10;

      		    if (~bfm_or_mon)
      		    begin //{

      		      lh_common_mon_trans.gen3_expected_c0_training_status[mon_type][lane_num] = 2'b10;

		      if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      begin //{
      		        current_c0_coeff_update_state = NOT_UPDATED;
		      end //}

      		    end //}
		    else
		    begin //{

		      if (~lh_trans.gen3_training_cmd_set[lane_num])
		      begin //{
      		        current_c0_coeff_update_state = NOT_UPDATED;
		      end //}

		    end //}

	    	  end //}

      endcase

      //if (prev_dme_train_state != current_dme_train_state && (current_dme_train_state == TRAINED || prev_dme_train_state == TRAINED))
      //  `uvm_info("SRIO_LANE_HANDLER : GEN3_DME_TRAIN_SM", $sformatf(" lane_trained[%0d] is %0d Next dme train state is %0s", lane_num, lh_trans.lane_trained[lane_num], current_dme_train_state.name()), UVM_LOW)

      if (~bfm_or_mon && prev_c0_coeff_update_state != current_c0_coeff_update_state)
        current_c0_coeff_update_state_q.push_back(current_c0_coeff_update_state);

    end //}

  end //}

endtask : gen3_c0_coeff_update_sm




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_cp1_coeff_update_sm
/// Description : This is the coefficient update state machine for tap CP1. The state machine
/// is defined in the 802.3-2008 specification.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_cp1_coeff_update_sm();

#1;
  if (~srio_if.srio_rst_n)
  begin //{

    current_cp1_coeff_update_state = NOT_UPDATED;

    if (bfm_or_mon)
    begin //{
      cp1_preset_value = lh_config.bfm_dme_training_cp1_preset_value;
      cp1_init_value = lh_config.bfm_dme_training_cp1_init_value;
      cp1_max_limit = lh_config.bfm_dme_training_cp1_max_value;
      cp1_min_limit = lh_config.bfm_dme_training_cp1_min_value;
    end //}
    else if (mon_type && lh_env_config.srio_tx_mon_if == DUT)
    begin //{
      cp1_preset_value = lh_config.bfm_dme_training_cp1_preset_value;
      cp1_init_value = lh_config.bfm_dme_training_cp1_init_value;
      cp1_max_limit = lh_config.bfm_dme_training_cp1_max_value;
      cp1_min_limit = lh_config.bfm_dme_training_cp1_min_value;
    end //}
    else if (mon_type && lh_env_config.srio_tx_mon_if == BFM)
    begin //{
      cp1_preset_value = lh_config.lp_dme_training_cp1_preset_value;
      cp1_init_value = lh_config.lp_dme_training_cp1_init_value;
      cp1_max_limit = lh_config.lp_dme_training_cp1_max_value;
      cp1_min_limit = lh_config.lp_dme_training_cp1_min_value;
    end //}
    else if (~mon_type && lh_env_config.srio_rx_mon_if == DUT)
    begin //{
      cp1_preset_value = lh_config.bfm_dme_training_cp1_preset_value;
      cp1_init_value = lh_config.bfm_dme_training_cp1_init_value;
      cp1_max_limit = lh_config.bfm_dme_training_cp1_max_value;
      cp1_min_limit = lh_config.bfm_dme_training_cp1_min_value;
    end //}
    else if (~mon_type && lh_env_config.srio_rx_mon_if == BFM)
    begin //{
      cp1_preset_value = lh_config.lp_dme_training_cp1_preset_value;
      cp1_init_value = lh_config.lp_dme_training_cp1_init_value;
      cp1_max_limit = lh_config.lp_dme_training_cp1_max_value;
      cp1_min_limit = lh_config.lp_dme_training_cp1_min_value;
    end //}

    if (~bfm_or_mon)
      current_cp1_coeff_update_state_q.push_back(current_cp1_coeff_update_state);

  end //}

  forever
  begin //{

    wait (lh_trans.frame_lock[lane_num] == 1);

    @(negedge dme_frame_divide_clk or negedge srio_if.srio_rst_n);

    if (~srio_if.srio_rst_n || lh_trans.mr_restart_training)
    begin //{

      prev_cp1_coeff_update_state = current_cp1_coeff_update_state;

      current_cp1_coeff_update_state = NOT_UPDATED;
      lh_trans.gen3_cp1_coeff_status[lane_num] = 2'b00;

      if (~bfm_or_mon)
      begin //{
        lh_common_mon_trans.gen3_expected_cp1_training_status[~mon_type][lane_num] = 2'b00;
      end //}

      if (~bfm_or_mon && prev_cp1_coeff_update_state != current_cp1_coeff_update_state)
        current_cp1_coeff_update_state_q.push_back(current_cp1_coeff_update_state);

    end //}
    else
    begin //{

      //`uvm_info("SRIO_LANE_HANDLER : GEN3_CW_TRAIN_SM", $sformatf(" lane_trained[%0d] is %0d Present cw train state is %0s", lane_num, lh_trans.lane_trained[lane_num], current_dme_train_state.name()), UVM_LOW)

      prev_cp1_coeff_update_state = current_cp1_coeff_update_state;

      case (current_cp1_coeff_update_state)

	NOT_UPDATED : begin //{

      			lh_trans.gen3_cp1_coeff_status[lane_num] = 2'b00;

      			if (~bfm_or_mon)
      			begin //{

      			  lh_common_mon_trans.gen3_expected_cp1_training_status[mon_type][lane_num] = 2'b00;

		      	  if (lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      	  begin //{
      		      	    current_cp1_coeff_update_state = UPDATE_COEFF;
		      	  end //}

      			end //}
			else
			begin //{

		      	  if (lh_trans.gen3_training_cmd_set[lane_num])
		      	  begin //{
      		      	    current_cp1_coeff_update_state = UPDATE_COEFF;
		      	  end //}

			end //}

		      end //}

	UPDATE_COEFF : begin //{

      			if (~bfm_or_mon)
      			begin //{

		      	  if (lh_common_mon_trans.gen3_c0_training_cmd[~mon_type][lane_num] == 3'b110)	// preset
		      	  begin //{
      		      	    new_cp1_coeff = cp1_preset_value;
		      	  end //}
		      	  else if (lh_common_mon_trans.gen3_c0_training_cmd[~mon_type][lane_num] == 3'b101) // Initialize
		      	  begin //{
      		      	    new_cp1_coeff = cp1_init_value;
		      	  end //}
		      	  else if (lh_common_mon_trans.gen3_cp1_training_cmd[~mon_type][lane_num] == 2'b10) // Increment
		      	  begin //{
      		      	    new_cp1_coeff = (new_cp1_coeff < cp1_max_limit) ? new_cp1_coeff+1 : cp1_max_limit;
		      	  end //}
		      	  else if (lh_common_mon_trans.gen3_cp1_training_cmd[~mon_type][lane_num] == 2'b01) // decrement
		      	  begin //{
      		      	    new_cp1_coeff = (new_cp1_coeff > cp1_min_limit) ? new_cp1_coeff-1 : cp1_min_limit;
		      	  end //}

      			end //}
			else
			begin //{


		      	  if (lh_trans.gen3_training_equalizer_cmd[lane_num] == 3'b110)	// preset
		      	  begin //{
      		      	    new_cp1_coeff = cp1_preset_value;
		      	  end //}
		      	  else if (lh_trans.gen3_training_equalizer_cmd[lane_num] == 3'b101) // Initialize
		      	  begin //{
      		      	    new_cp1_coeff = cp1_init_value;
		      	  end //}
		      	  else if (lh_trans.gen3_training_equalizer_cp1_cmd[lane_num] == 2'b10) // Increment
		      	  begin //{
      		      	    new_cp1_coeff = (new_cp1_coeff < cp1_max_limit) ? new_cp1_coeff+1 : cp1_max_limit;
		      	  end //}
		      	  else if (lh_trans.gen3_training_equalizer_cp1_cmd[lane_num] == 2'b01) // decrement
		      	  begin //{
      		      	    new_cp1_coeff = (new_cp1_coeff > cp1_min_limit) ? new_cp1_coeff-1 : cp1_min_limit;
		      	  end //}

			end //}

			if (new_cp1_coeff >= cp1_max_limit)
			  current_cp1_coeff_update_state = MAXIMUM;
			else if ((new_cp1_coeff > cp1_min_limit) && (new_cp1_coeff < cp1_max_limit))
			  current_cp1_coeff_update_state = UPDATED;
			else if (new_cp1_coeff <= cp1_max_limit)
			  current_cp1_coeff_update_state = MINIMUM;

		      end //}

	MAXIMUM : begin //{

      		    lh_trans.gen3_cp1_coeff_status[lane_num] = 2'b11;

      		    if (~bfm_or_mon)
      		    begin //{

      		      lh_common_mon_trans.gen3_expected_cp1_training_status[mon_type][lane_num] = 2'b11;

		      if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      begin //{
      		        current_cp1_coeff_update_state = NOT_UPDATED;
		      end //}

      		    end //}
		    else
		    begin //{

		      if (~lh_trans.gen3_training_cmd_set[lane_num])
		      begin //{
      		        current_cp1_coeff_update_state = NOT_UPDATED;
		      end //}

		    end //}

	    	  end //}

	UPDATED : begin //{

      		    lh_trans.gen3_cp1_coeff_status[lane_num] = 2'b01;

      		    if (~bfm_or_mon)
      		    begin //{

      		      lh_common_mon_trans.gen3_expected_cp1_training_status[mon_type][lane_num] = 2'b01;

		      if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      begin //{
      		        current_cp1_coeff_update_state = NOT_UPDATED;
		      end //}

      		    end //}
		    else
		    begin //{

		      if (~lh_trans.gen3_training_cmd_set[lane_num])
		      begin //{
      		        current_cp1_coeff_update_state = NOT_UPDATED;
		      end //}

		    end //}

	    	  end //}

	MINIMUM : begin //{

      		    lh_trans.gen3_cp1_coeff_status[lane_num] = 2'b10;

      		    if (~bfm_or_mon)
      		    begin //{

      		      lh_common_mon_trans.gen3_expected_cp1_training_status[mon_type][lane_num] = 2'b10;

		      if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      begin //{
      		        current_cp1_coeff_update_state = NOT_UPDATED;
		      end //}

      		    end //}
		    else
		    begin //{

		      if (~lh_trans.gen3_training_cmd_set[lane_num])
		      begin //{
      		        current_cp1_coeff_update_state = NOT_UPDATED;
		      end //}

		    end //}

	    	  end //}

      endcase

      //if (prev_dme_train_state != current_dme_train_state && (current_dme_train_state == TRAINED || prev_dme_train_state == TRAINED))
      //  `uvm_info("SRIO_LANE_HANDLER : GEN3_DME_TRAIN_SM", $sformatf(" lane_trained[%0d] is %0d Next dme train state is %0s", lane_num, lh_trans.lane_trained[lane_num], current_dme_train_state.name()), UVM_LOW)

      if (~bfm_or_mon && prev_cp1_coeff_update_state != current_cp1_coeff_update_state)
        current_cp1_coeff_update_state_q.push_back(current_cp1_coeff_update_state);


    end //}

  end //}

endtask : gen3_cp1_coeff_update_sm




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_cn1_coeff_update_sm
/// Description : This is the coefficient update state machine for tap CN1. The state machine
/// is defined in the 802.3-2008 specification.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_cn1_coeff_update_sm();

#1;
  if (~srio_if.srio_rst_n)
  begin //{

    current_cn1_coeff_update_state = NOT_UPDATED;

    if (bfm_or_mon)
    begin //{
      cn1_preset_value = lh_config.bfm_dme_training_cn1_preset_value;
      cn1_init_value = lh_config.bfm_dme_training_cn1_init_value;
      cn1_max_limit = lh_config.bfm_dme_training_cn1_max_value;
      cn1_min_limit = lh_config.bfm_dme_training_cn1_min_value;
    end //}
    else if (mon_type && lh_env_config.srio_tx_mon_if == DUT)
    begin //{
      cn1_preset_value = lh_config.bfm_dme_training_cn1_preset_value;
      cn1_init_value = lh_config.bfm_dme_training_cn1_init_value;
      cn1_max_limit = lh_config.bfm_dme_training_cn1_max_value;
      cn1_min_limit = lh_config.bfm_dme_training_cn1_min_value;
    end //}
    else if (mon_type && lh_env_config.srio_tx_mon_if == BFM)
    begin //{
      cn1_preset_value = lh_config.lp_dme_training_cn1_preset_value;
      cn1_init_value = lh_config.lp_dme_training_cn1_init_value;
      cn1_max_limit = lh_config.lp_dme_training_cn1_max_value;
      cn1_min_limit = lh_config.lp_dme_training_cn1_min_value;
    end //}
    else if (~mon_type && lh_env_config.srio_rx_mon_if == DUT)
    begin //{
      cn1_preset_value = lh_config.bfm_dme_training_cn1_preset_value;
      cn1_init_value = lh_config.bfm_dme_training_cn1_init_value;
      cn1_max_limit = lh_config.bfm_dme_training_cn1_max_value;
      cn1_min_limit = lh_config.bfm_dme_training_cn1_min_value;
    end //}
    else if (~mon_type && lh_env_config.srio_rx_mon_if == BFM)
    begin //{
      cn1_preset_value = lh_config.lp_dme_training_cn1_preset_value;
      cn1_init_value = lh_config.lp_dme_training_cn1_init_value;
      cn1_max_limit = lh_config.lp_dme_training_cn1_max_value;
      cn1_min_limit = lh_config.lp_dme_training_cn1_min_value;
    end //}

    if (~bfm_or_mon)
      current_cn1_coeff_update_state_q.push_back(current_cn1_coeff_update_state);

  end //}

  forever
  begin //{

    wait (lh_trans.frame_lock[lane_num] == 1);

    @(negedge dme_frame_divide_clk or negedge srio_if.srio_rst_n);

    if (~srio_if.srio_rst_n || lh_trans.mr_restart_training)
    begin //{

      prev_cn1_coeff_update_state = current_cn1_coeff_update_state;

      current_cn1_coeff_update_state = NOT_UPDATED;
      lh_trans.gen3_cn1_coeff_status[lane_num] = 2'b00;

      if (~bfm_or_mon)
      begin //{
        lh_common_mon_trans.gen3_expected_cn1_training_status[~mon_type][lane_num] = 2'b00;
      end //}

      if (~bfm_or_mon && prev_cn1_coeff_update_state != current_cn1_coeff_update_state)
        current_cn1_coeff_update_state_q.push_back(current_cn1_coeff_update_state);

    end //}
    else
    begin //{

      //`uvm_info("SRIO_LANE_HANDLER : GEN3_CW_TRAIN_SM", $sformatf(" lane_trained[%0d] is %0d Present cw train state is %0s", lane_num, lh_trans.lane_trained[lane_num], current_dme_train_state.name()), UVM_LOW)

      prev_cn1_coeff_update_state = current_cn1_coeff_update_state;

      case (current_cn1_coeff_update_state)

	NOT_UPDATED : begin //{

      			lh_trans.gen3_cn1_coeff_status[lane_num] = 2'b00;

      			if (~bfm_or_mon)
      			begin //{

      			  lh_common_mon_trans.gen3_expected_cn1_training_status[mon_type][lane_num] = 2'b00;

		      	  if (lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      	  begin //{
      		      	    current_cn1_coeff_update_state = UPDATE_COEFF;
		      	  end //}

      			end //}
			else
			begin //{

		      	  if (lh_trans.gen3_training_cmd_set[lane_num])
		      	  begin //{
      		      	    current_cn1_coeff_update_state = UPDATE_COEFF;
		      	  end //}

			end //}

		      end //}

	UPDATE_COEFF : begin //{

      			if (~bfm_or_mon)
      			begin //{

		      	  if (lh_common_mon_trans.gen3_c0_training_cmd[~mon_type][lane_num] == 3'b110)	// preset
		      	  begin //{
      		      	    new_cn1_coeff = cn1_preset_value;
		      	  end //}
		      	  else if (lh_common_mon_trans.gen3_c0_training_cmd[~mon_type][lane_num] == 3'b101) // Initialize
		      	  begin //{
      		      	    new_cn1_coeff = cn1_init_value;
		      	  end //}
		      	  else if (lh_common_mon_trans.gen3_cn1_training_cmd[~mon_type][lane_num] == 2'b10) // Increment
		      	  begin //{
      		      	    new_cn1_coeff = (new_cn1_coeff < cn1_max_limit) ? new_cn1_coeff+1 : cn1_max_limit;
		      	  end //}
		      	  else if (lh_common_mon_trans.gen3_cn1_training_cmd[~mon_type][lane_num] == 2'b01) // decrement
		      	  begin //{
      		      	    new_cn1_coeff = (new_cn1_coeff > cn1_min_limit) ? new_cn1_coeff-1 : cn1_min_limit;
		      	  end //}

      			end //}
			else
			begin //{


		      	  if (lh_trans.gen3_training_equalizer_cmd[lane_num] == 3'b110)	// preset
		      	  begin //{
      		      	    new_cn1_coeff = cn1_preset_value;
		      	  end //}
		      	  else if (lh_trans.gen3_training_equalizer_cmd[lane_num] == 3'b101) // Initialize
		      	  begin //{
      		      	    new_cn1_coeff = cn1_init_value;
		      	  end //}
		      	  else if (lh_trans.gen3_training_equalizer_cn1_cmd[lane_num] == 2'b10) // Increment
		      	  begin //{
      		      	    new_cn1_coeff = (new_cn1_coeff < cn1_max_limit) ? new_cn1_coeff+1 : cn1_max_limit;
		      	  end //}
		      	  else if (lh_trans.gen3_training_equalizer_cn1_cmd[lane_num] == 2'b01) // decrement
		      	  begin //{
      		      	    new_cn1_coeff = (new_cn1_coeff > cn1_min_limit) ? new_cn1_coeff-1 : cn1_min_limit;
		      	  end //}

			end //}

			if (new_cn1_coeff >= cn1_max_limit)
			  current_cn1_coeff_update_state = MAXIMUM;
			else if ((new_cn1_coeff > cn1_min_limit) && (new_cn1_coeff < cn1_max_limit))
			  current_cn1_coeff_update_state = UPDATED;
			else if (new_cn1_coeff <= cn1_max_limit)
			  current_cn1_coeff_update_state = MINIMUM;

		      end //}

	MAXIMUM : begin //{

      		    lh_trans.gen3_cn1_coeff_status[lane_num] = 2'b11;

      		    if (~bfm_or_mon)
      		    begin //{

      		      lh_common_mon_trans.gen3_expected_cn1_training_status[mon_type][lane_num] = 2'b11;

		      if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      begin //{
      		        current_cn1_coeff_update_state = NOT_UPDATED;
		      end //}

      		    end //}
		    else
		    begin //{

		      if (~lh_trans.gen3_training_cmd_set[lane_num])
		      begin //{
      		        current_cn1_coeff_update_state = NOT_UPDATED;
		      end //}

		    end //}

	    	  end //}

	UPDATED : begin //{

      		    lh_trans.gen3_cn1_coeff_status[lane_num] = 2'b01;

      		    if (~bfm_or_mon)
      		    begin //{

      		      lh_common_mon_trans.gen3_expected_cn1_training_status[mon_type][lane_num] = 2'b01;

		      if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      begin //{
      		        current_cn1_coeff_update_state = NOT_UPDATED;
		      end //}

      		    end //}
		    else
		    begin //{

		      if (~lh_trans.gen3_training_cmd_set[lane_num])
		      begin //{
      		        current_cn1_coeff_update_state = NOT_UPDATED;
		      end //}

		    end //}

	    	  end //}

	MINIMUM : begin //{

      		    lh_trans.gen3_cn1_coeff_status[lane_num] = 2'b10;

      		    if (~bfm_or_mon)
      		    begin //{

      		      lh_common_mon_trans.gen3_expected_cn1_training_status[mon_type][lane_num] = 2'b10;

		      if (~lh_common_mon_trans.gen3_training_cmd_outstanding[~mon_type][lane_num])
		      begin //{
      		        current_cn1_coeff_update_state = NOT_UPDATED;
		      end //}

      		    end //}
		    else
		    begin //{

		      if (~lh_trans.gen3_training_cmd_set[lane_num])
		      begin //{
      		        current_cn1_coeff_update_state = NOT_UPDATED;
		      end //}

		    end //}

	    	  end //}

      endcase

      //if (prev_dme_train_state != current_dme_train_state && (current_dme_train_state == TRAINED || prev_dme_train_state == TRAINED))
      //  `uvm_info("SRIO_LANE_HANDLER : GEN3_DME_TRAIN_SM", $sformatf(" lane_trained[%0d] is %0d Next dme train state is %0s", lane_num, lh_trans.lane_trained[lane_num], current_dme_train_state.name()), UVM_LOW)

      if (~bfm_or_mon && prev_cn1_coeff_update_state != current_cn1_coeff_update_state)
        current_cn1_coeff_update_state_q.push_back(current_cn1_coeff_update_state);

    end //}

  end //}

endtask : gen3_cn1_coeff_update_sm




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : cw_lock_sm
/// Description : Implements the codeword lock state machine as defined in the GEN3.0 specification
/// Waiting for the next negedge of clk or reset is bypassed when intermediate states are encountered
/// by the state machine.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::cw_lock_sm();

  //int CW_counter;
  //int V_counter;
  //int IV_counter;

#1;
  if (~srio_if.srio_rst_n)
  begin //{
    current_cw_lock_state = NO_LOCK;
    if (~bfm_or_mon)
      current_cw_lock_state_q.push_back(current_cw_lock_state);
    // questasim and vcs doesn't work properly on associatuve array methods
    // Hence, a work-around is done here by setting the array values to 1 and
    // then clearing it immediately.
    lh_trans.cw_lock[lane_num] = 1;
    lh_trans.cw_lock[lane_num] = 0;

    lh_trans.rcvr_trained[lane_num] = 1;
    if (lh_config.aet_en)
      lh_trans.rcvr_trained[lane_num] = 0;

    lh_trans.signal_detect[lane_num] = 1;
    lh_trans.signal_detect[lane_num] = 0;
    lh_trans.lane_ready[lane_num] = 1;
    lh_trans.lane_ready[lane_num] = 0;
    CW_counter = 0;
    V_counter = 0;
  end //}

  forever
  begin //{

    // In the following conditions, there's no need to wait for the negedge of clock, 
    // as it would lead to missing of alternate data
    if (!(prev_cw_lock_state == NO_LOCK_1 && current_cw_lock_state == NO_LOCK_2) && !(prev_cw_lock_state == LOCK && current_cw_lock_state == LOCK_1) && !(prev_cw_lock_state == LOCK_2 && current_cw_lock_state == LOCK_1) && !(prev_cw_lock_state == LOCK_3 && current_cw_lock_state == LOCK_1))
      @(negedge divide_clk or negedge srio_if.srio_rst_n or negedge lh_trans.signal_detect[lane_num] or posedge lh_trans.force_no_lock[lane_num]);

    if (~srio_if.srio_rst_n || ~lh_trans.signal_detect[lane_num] || lh_trans.force_no_lock[lane_num])
    begin //{

      prev_cw_lock_state = current_cw_lock_state;

      current_cw_lock_state = NO_LOCK;
      lh_trans.cw_lock[lane_num] = 0;
      CW_counter = 0;
      V_counter = 0;
      IV_counter = 0;
      s2p_lock = 0;

      if (~bfm_or_mon)
      begin //{
        if (lh_common_mon_trans.sc_os_cnt[~mon_type] > 0 && lh_common_mon_trans.sc_os_cnt[~mon_type] < 8)
        begin //{
          `uvm_warning("SRIO_PL_LANE_HANDLER : SC_OS_AFTER_PORT_ENTERING_SILENCE", $sformatf(" Spec reference 5.8.2. Atleast 8 Status-Control ordered sequence has to be transmitted with port/lane entering silence set before entering into SILENT state.. No of Status-Control ordererd sequence sent with port/lane entering silence field set is %0d", lh_common_mon_trans.sc_os_cnt[~mon_type]))
        end //}
        lh_common_mon_trans.sc_os_cnt[~mon_type] = 0;
      end //}
      if (~bfm_or_mon && prev_cw_lock_state != current_cw_lock_state)
	current_cw_lock_state_q.push_back(current_cw_lock_state);

    end //}
    else
    begin //{

      //`uvm_info("SRIO_LANE_HANDLER : LOCK_SM", $sformatf(" cw_lock[%0d] is %0d Present lock state is %0s", lane_num, lh_trans.cw_lock[lane_num], current_cw_lock_state.name()), UVM_LOW)

      prev_cw_lock_state = current_cw_lock_state;

      case (current_cw_lock_state)

	NO_LOCK : begin //{

		   //$display($time, " : Entered NO_LOCK in lane_num %0d", lane_num);

		     lh_trans.cw_lock[lane_num] = 0;

		     current_cw_lock_state = NO_LOCK_1;
		     if (~bfm_or_mon)
		     begin //{
		       if (lh_common_mon_trans.sc_os_cnt[~mon_type] > 0 && lh_common_mon_trans.sc_os_cnt[~mon_type] < 8)
		       begin //{
		         `uvm_warning("SRIO_PL_LANE_HANDLER : SC_OS_AFTER_PORT_ENTERING_SILENCE", $sformatf(" Spec reference 5.8.2. Atleast 8 Status-Control ordered sequence has to be transmitted with port/lane entering silence set before entering into SILENT state.. No of Status-Control ordererd sequence sent with port/lane entering silence field set is %0d", lh_common_mon_trans.sc_os_cnt[~mon_type]))
		       end //}
		       lh_common_mon_trans.sc_os_cnt[~mon_type] = 0;
		     end //}

		   end //}

	NO_LOCK_1 : begin //{

		      lh_trans.cw_lock[lane_num] = 0;
      		      V_counter = 0;

		      current_cw_lock_state = NO_LOCK_2;

		    end //}

	NO_LOCK_2 : begin //{

		      lh_trans.cw_lock[lane_num] = 0;

		      if (lane_data_ins.brc3_cg[1] == ~lane_data_ins.brc3_cg[2])
			current_cw_lock_state = NO_LOCK_3;
		      else
                       begin//{
			current_cw_lock_state = SLIP_ALIGNMENT;
                        if(lh_config.parallel_cw_slip_adj_en && lh_env_config.srio_interface_mode == SRIO_PARALLEL)
                         begin//{
                          note_bit_3=67;
                          for(int k=0;k<=note_bit_3;k++)
                           begin//{
	                    if (sixty_seven_bit_data[1] == ~sixty_seven_bit_data[2])
                             begin//{
	                      s2p_lock = 1;
                              note_bit_1=note_bit_1+k;
                              if(k==67)
                               note_bit_1=note_bit_1;
                              if(note_bit_1>67) 
                               note_bit_1=note_bit_1-67;
                              break;
                             end//}
                            else
                             begin//{
                              if(k!=67)
                               begin//{
                                sixty_seven_bit_data=sixty_seven_bit_data<<1;
                                sixty_seven_bit_data[66]=sixty_seven_bit_data_tmp[0];
                                sixty_seven_bit_data_tmp=sixty_seven_bit_data_tmp<<1;
                               end//}
                             end//}
                           end//}
                         if(s2p_lock)
	                    	current_cw_lock_state = NO_LOCK_3;
                         else
	                    	current_cw_lock_state = SLIP_ALIGNMENT;
                       end//}
                      end//}

		    end //}

	NO_LOCK_3 : begin //{

		      lh_trans.cw_lock[lane_num] = 0;
      		      V_counter++;

		      if (V_counter < lh_config.brc3_v_cnt_threshold)
		        current_cw_lock_state = NO_LOCK_2;
		      else
		        current_cw_lock_state = LOCK;

		    end //}

	LOCK : begin //{

		   //$display($time, " : Entered LOCK in lane_num %0d", lane_num);

	         lh_trans.cw_lock[lane_num] = 1;
      	         CW_counter = 0;
      	         IV_counter = 0;

	         current_cw_lock_state = LOCK_1;

	       end //}

	LOCK_1 : begin //{

		   //$display($time, " : Entered LOCK_1 in lane_num %0d", lane_num);

	           lh_trans.cw_lock[lane_num] = 1;

		   if (lane_data_ins.brc3_cg[1] == ~lane_data_ins.brc3_cg[2])
		     current_cw_lock_state = LOCK_3;
		   else
		     current_cw_lock_state = LOCK_2;

	       	 end //}

	LOCK_2 : begin //{

		   //$display($time, " : Entered LOCK_2 in lane_num %0d", lane_num);

	           lh_trans.cw_lock[lane_num] = 1;
      	           CW_counter++;
      	           IV_counter++;


		   if (IV_counter < lh_config.lock_break_threshold)
	             current_cw_lock_state = LOCK_1;
		   else
	             current_cw_lock_state = NO_LOCK;

	       	 end //}

	LOCK_3 : begin //{

		   //$display($time, " : Entered LOCK_3 in lane_num %0d", lane_num);

	           lh_trans.cw_lock[lane_num] = 1;
      	           CW_counter++;

		   if (CW_counter < lh_config.brc3_v_cnt_threshold)
	             current_cw_lock_state = LOCK_1;
		   else
	             current_cw_lock_state = LOCK;

	       	 end //}

	SLIP_ALIGNMENT : begin //{

		   	   //$display($time, " : Entered SLIP_ALIGNMENT in lane_num %0d", lane_num);

			   s2p_lock = 0;

	           	   current_cw_lock_state = NO_LOCK_1;

	       	 	 end //}

      endcase

      //if (prev_cw_lock_state != current_cw_lock_state && (current_cw_lock_state == LOCK || prev_cw_lock_state == LOCK))
      //  `uvm_info("SRIO_LANE_HANDLER : LOCK_SM", $sformatf(" cw_lock[%0d] is %0d Next lock state is %0s", lane_num, lh_trans.cw_lock[lane_num], current_cw_lock_state.name()), UVM_LOW)

      if (~bfm_or_mon && prev_cw_lock_state != current_cw_lock_state)
	current_cw_lock_state_q.push_back(current_cw_lock_state);

    end //}

  end //}

endtask : cw_lock_sm



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_lane_sync_sm
/// Description : Implements the lane sync state machine for GEN3.0 device.
/// Waiting for the next negedge of clk or reset is bypassed when intermediate states are encountered
/// by the state machine.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_lane_sync_sm();

  int DS_counter;

#1;
  if (~srio_if.srio_rst_n)
  begin //{
    current_sync_state = NO_SYNC;
    if (~bfm_or_mon)
      current_sync_state_q.push_back(current_sync_state);
    // questasim and vcs doesn't work properly on associatuve array methods
    // Hence, a work-around is done here by setting the array values to 1 and
    // then clearing it immediately.
    lh_trans.lane_sync[lane_num] = 1;
    lh_trans.lane_sync[lane_num] = 0;

    lh_trans.force_no_lock[lane_num] = 1;
    lh_trans.force_no_lock[lane_num] = 0;

    lh_trans.frame_lock[lane_num] = 1;
    lh_trans.frame_lock[lane_num] = 0;

    DS_counter = 0;

  end //}

  if (~bfm_or_mon)
    update_ls0_lane_num_field();

  forever
  begin //{

    // In the following conditions, there's no need to wait for the negedge of clock, 
    // as it would lead to missing of alternate data
    if (!(prev_sync_state == NO_SYNC_1 && current_sync_state == NO_SYNC_2) && !(prev_sync_state == NO_SYNC_3 && current_sync_state == NO_SYNC_2) && !(prev_sync_state == NO_SYNC_4 && current_sync_state == NO_SYNC_2))
      @(negedge divide_clk or negedge srio_if.srio_rst_n or negedge lh_trans.cw_lock[lane_num]);

    if (~srio_if.srio_rst_n || ~lh_trans.cw_lock[lane_num])
    begin //{

      prev_sync_state = current_sync_state;

      current_sync_state = NO_SYNC;
      lh_trans.lane_sync[lane_num] = 0;
      lh_trans.force_no_lock[lane_num] = 0;
      DS_counter = 0;

      if (~bfm_or_mon && prev_sync_state != current_sync_state)
	current_sync_state_q.push_back(current_sync_state);

    end //}
    else
    begin //{

      //`uvm_info("SRIO_LANE_HANDLER : SYNC_SM", $sformatf(" lane_sync[%0d] is %0d Present sync state is %0s", lane_num, lh_trans.lane_sync[lane_num], current_sync_state.name()), UVM_LOW)

      prev_sync_state = current_sync_state;

      case (current_sync_state)

	NO_SYNC : begin //{

		   //$display($time, " : Entered NO_SYNC in lane_num %0d", lane_num);

		     lh_trans.lane_sync[lane_num] = 0;
		     lh_trans.force_no_lock[lane_num] = 0;

		     if (lh_trans.cw_lock[lane_num])
		       current_sync_state = NO_SYNC_1;

		   end //}

	NO_SYNC_1 : begin //{

		      lh_trans.lane_sync[lane_num] = 0;
      		      DS_counter = 0;

		      current_sync_state = NO_SYNC_2;

		    end //}

	NO_SYNC_2 : begin //{

		      lh_trans.lane_sync[lane_num] = 0;

		      current_sync_state = NO_SYNC_3;

		    end //}

	NO_SYNC_3 : begin //{

		      lh_trans.lane_sync[lane_num] = 0;

		      if (sync_sm_descr_sync)
		        current_sync_state = NO_SYNC_4;
		      else if (sync_sm_descr_err)
		        current_sync_state = NO_SYNC_1;
		      else
		        current_sync_state = NO_SYNC_2;

		    end //}

	NO_SYNC_4 : begin //{

		      lh_trans.lane_sync[lane_num] = 0;
		      DS_counter++;

		      if (DS_counter < lh_config.brc3_ds_cnt_threshold)
		        current_sync_state = NO_SYNC_2;
		      else
		        current_sync_state = SYNC;

		    end //}

	SYNC : begin //{

	         lh_trans.lane_sync[lane_num] = 1;

		 if (lh_trans.from_sc_port_silence || lh_trans.from_sc_lane_silence[lane_num])
	           current_sync_state = SYNC_1;

	       end //}

	SYNC_1 : begin //{

		   //$display($time, " : Entered SYNC_1 in lane_num %0d", lane_num);

	           lh_trans.lane_sync[lane_num] = 1;
		   sync1_state_ui_cnt++;

		   if (sync1_state_ui_cnt == lh_config.sync1_state_ui_cnt_threshold)
		   begin //{
		     sync1_state_ui_cnt = 0;
	             current_sync_state = SYNC_2;
		   end //}

	       	 end //}

	SYNC_2 : begin //{

		   //$display($time, " : Entered SYNC_2 in lane_num %0d", lane_num);

	           lh_trans.lane_sync[lane_num] = 1;
	           lh_trans.force_no_lock[lane_num] = 1;

	       	 end //}

      endcase

      if (prev_sync_state != current_sync_state && (current_sync_state == SYNC || prev_sync_state == SYNC))
        `uvm_info("SRIO_LANE_HANDLER : SYNC_SM", $sformatf(" lane_sync[%0d] is %0d Next sync state is %0s", lane_num, lh_trans.lane_sync[lane_num], current_sync_state.name()), UVM_LOW)

      if (~bfm_or_mon && prev_sync_state != current_sync_state)
	current_sync_state_q.push_back(current_sync_state);

    end //}

   // if (lh_trans.lane_sync[lane_num] == 1)
      temp_lane_data_ins = new lane_data_ins;
      //$cast(temp_lane_data_ins, lane_data_ins.clone());
      srio_rx_lane_event.trigger(temp_lane_data_ins);
//	if (~bfm_or_mon && ~mon_type)
//	$display($time, " lane_num is %0d, mon_type is %0d. Event triggered from sync sm. lane_data_ins.character is %0h temp_lane_data_ins.character is %0h", lane_num, mon_type, lane_data_ins.character, temp_lane_data_ins.character);

  end //}

endtask : gen3_lane_sync_sm



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_cw_training_sm
/// Description : Implements the CW training / short-run training state machine for GEN3.0 device.
/// Since the complete CW training logic is also available as a part of long-run training state 
/// machine, the below method is used for both short-run training as well as for CW training part of
/// long-run training. The switching is done such that,if long-run mode is active and if the long-run
/// training state reaches either CW_TRAINING_0 state or TRAINED state, this method will become active.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_cw_training_sm();

#1;
  if (~srio_if.srio_rst_n)
  begin //{
    current_cw_train_state = UNTRAINED;

    if (~bfm_or_mon)
      current_cw_train_state_q.push_back(current_cw_train_state);

    // questasim and vcs doesn't work properly on associatuve array methods
    // Hence, a work-around is done here by setting the array values to 1 and
    // then clearing it immediately.
    lh_trans.lane_retraining[lane_num] = 1;
    lh_trans.lane_retraining[lane_num] = 0;

    lh_trans.lane_trained[lane_num] = 1;
    lh_trans.lane_trained[lane_num] = 0;

    lh_trans.from_sc_lane_trained[lane_num] = 1;
    lh_trans.from_sc_lane_trained[lane_num] = 0;

    lh_trans.from_sc_lane_silence[lane_num] = 1;
    lh_trans.from_sc_lane_silence[lane_num] = 0;

    lh_trans.gen3_training_equalizer_tap[lane_num] = 1;
    lh_trans.gen3_training_equalizer_cmd[lane_num] = 1;
    lh_trans.gen3_training_equalizer_status[lane_num] = 1;

    lh_trans.dme_mode[lane_num] = 1;
    lh_trans.train_lane[lane_num] = 1;
    lh_trans.retrain_lane[lane_num] = 1;
    lh_trans.train_timer_en[lane_num] = 1;
    lh_trans.train_timer_done[lane_num] = 1;

    lh_trans.force_drvr_oe [lane_num] = 1;
    lh_trans.drvr_oe [lane_num] = 1;

    lh_trans.keep_alive [lane_num] = 1;

    lh_trans.lane_degraded [lane_num] = 1;
    lh_trans.retrain_fail [lane_num] = 1;
    lh_trans.training_fail [lane_num] = 1;

    lh_trans.gen3_training_equalizer_tap[lane_num] = 0;
    lh_trans.gen3_training_equalizer_cmd[lane_num] = 0;
    lh_trans.gen3_training_equalizer_status[lane_num] = 0;

    if (~lh_config.brc3_training_mode)
      lh_trans.dme_mode[lane_num] = 0;

    lh_trans.train_lane[lane_num] = 0;
    lh_trans.retrain_lane[lane_num] = 0;
    lh_trans.train_timer_en[lane_num] = 0;
    lh_trans.train_timer_done[lane_num] = 0;

    lh_trans.force_drvr_oe [lane_num] = 0;
    //lh_trans.drvr_oe [lane_num] = 0;

    lh_trans.keep_alive [lane_num] = 0;

    lh_trans.lane_degraded [lane_num] = 0;
    lh_trans.retrain_fail [lane_num] = 0;
    lh_trans.training_fail [lane_num] = 0;

    if (~bfm_or_mon)
    begin //{

      lh_common_mon_trans.gen3_training_cmd_outstanding[mon_type][lane_num] = 1;
      lh_common_mon_trans.gen3_training_status_received[mon_type][lane_num] = 1;
      lh_common_mon_trans.gen3_cmd_deassertion_timer_started[mon_type][lane_num] = 1;

      lh_common_mon_trans.gen3_training_cmd_outstanding[mon_type][lane_num] = 0;
      lh_common_mon_trans.gen3_training_status_received[mon_type][lane_num] = 0;
      lh_common_mon_trans.gen3_cmd_deassertion_timer_started[mon_type][lane_num] = 0;

    end //}

  end //}

  forever
  begin //{

    if (lh_config.brc3_training_mode && current_dme_train_state != CW_TRAINING_0 && current_dme_train_state != TRAINED)
    begin //{

      wait((~lh_trans.frame_lock[lane_num] && lh_trans.lane_sync[lane_num] && current_dme_train_state == CW_TRAINING_0) || (lh_trans.frame_lock[lane_num] && current_dme_train_state == TRAINED));
      current_cw_train_state = current_dme_train_state;

      if (~bfm_or_mon && prev_cw_train_state != current_cw_train_state)
	current_cw_train_state_q.push_back(current_cw_train_state);

    end //}

    @(negedge divide_clk or negedge srio_if.srio_rst_n);

    if (~srio_if.srio_rst_n || (lh_trans.current_init_state == SILENT))
    begin //{

      prev_cw_train_state = current_cw_train_state;

      current_cw_train_state = UNTRAINED;

      if (~bfm_or_mon && prev_cw_train_state != current_cw_train_state)
	current_cw_train_state_q.push_back(current_cw_train_state);

      if (~bfm_or_mon)
	update_ls1_idle3_training_type(3'b000);

      lh_trans.lane_trained[lane_num] = 0;

      lh_trans.force_drvr_oe[lane_num] = 0;

      if (~lh_config.brc3_training_mode)
        lh_trans.dme_mode[lane_num] = 0;

      lh_trans.train_lane[lane_num] = 0;
      lh_trans.retrain_lane[lane_num] = 0;
      lh_trans.train_timer_en[lane_num] = 0;

    end //}
    else
    begin //{

      //`uvm_info("SRIO_LANE_HANDLER : GEN3_CW_TRAIN_SM", $sformatf(" lane_trained[%0d] is %0d Present cw train state is %0s", lane_num, lh_trans.lane_trained[lane_num], current_cw_train_state.name()), UVM_LOW)

      prev_cw_train_state = current_cw_train_state;

      case (current_cw_train_state)

	UNTRAINED : begin //{

      		      lh_trans.force_drvr_oe[lane_num] = 0;
      		      lh_trans.train_lane[lane_num] = 0;
      		      lh_trans.retrain_lane[lane_num] = 0;
      		      lh_trans.train_timer_en[lane_num] = 0;

      		      if (~lh_config.brc3_training_mode)
      		      begin //{
      		        lh_trans.dme_mode[lane_num] = 0;
		        lh_trans.xmt_equalizer = "SR_initialize";
      		      end //}

		      if (lh_trans.drvr_oe[lane_num] & lh_trans.lane_sync[lane_num])
		      begin //{
      			current_cw_train_state = CW_TRAINING_0;
		      end //}

		      if (~bfm_or_mon)
			update_ls1_idle3_training_type(3'b000);

		    end //}

	CW_TRAINING_0 : begin //{

		      	  lh_trans.train_timer_en[lane_num] = 1;
      		      	  lh_trans.dme_mode[lane_num] = 0;

		      	  lh_trans.xmt_equalizer = "SR_initialize";

		      	  if (lh_trans.train_timer_done[lane_num])
		      	    current_cw_train_state = CW_TRAINING_FAIL;
		      	  else if (!lh_trans.train_timer_done[lane_num] & !lh_trans.lane_trained[lane_num])
		      	    current_cw_train_state = CW_TRAINING_1;

		          if (~bfm_or_mon)
		    	    update_ls1_idle3_training_type(3'b010);

		    	end //}

	CW_TRAINING_1 : begin //{

      		      	  lh_trans.training_fail[lane_num] = 0;
		      	  lh_trans.train_lane[lane_num] = 1;

		      	  if (lh_trans.train_timer_done[lane_num])
		      	    current_cw_train_state = CW_TRAINING_FAIL;
		      	  else if (!lh_trans.train_timer_done[lane_num] & !lh_trans.drvr_oe[lane_num])
		      	    current_cw_train_state = UNTRAINED;
		      	  else if (!lh_trans.train_timer_done[lane_num] & lh_trans.drvr_oe[lane_num] & lh_trans.lane_sync[lane_num]
					& lh_trans.lane_trained[lane_num] & lh_trans.from_sc_lane_trained[lane_num])
		      	    current_cw_train_state = TRAINED;

		          if (~bfm_or_mon)
		          begin //{
		    	    update_ls1_idle3_training_type(3'b010);
			    //if (current_cw_train_state == TRAINED)
		    	    //  update_ls1_idle3_cw_training_completed();
		          end //}

		    	end //}

	CW_TRAINING_FAIL : begin //{

      		      	     lh_trans.training_fail[lane_num] = 1;
		      	     current_cw_train_state = UNTRAINED;

		             if (~bfm_or_mon)
		             begin //{
		    	       update_ls1_idle3_training_type(3'b010);
      		      	       update_ls1_idle3_cw_training_state();
		             end //}

		           end //}

	TRAINED : begin //{

      		      lh_trans.force_drvr_oe[lane_num] = 0;
      		      lh_trans.train_lane[lane_num] = 0;
      		      lh_trans.retrain_lane[lane_num] = 0;
      		      lh_trans.train_timer_en[lane_num] = 0;
                      lh_trans.dme_mode[lane_num] = 0;

		      if (lh_config.brc3_training_mode)
		      begin //{
			if (bfm_or_mon)
      		          lh_trans.dme_wait_timer_en[lane_num] = 0;
			else
      		          lh_common_mon_trans.dme_wait_timer_en[mon_type][lane_num] = 0;
		      end //}

		      if (lh_trans.retrain)
		        current_cw_train_state = RETRAINING_0;
		      else if (lh_trans.keep_alive[lane_num] & !lh_trans.retrain)
		        current_cw_train_state = KEEP_ALIVE;

		      if (~bfm_or_mon)
		        update_ls1_idle3_training_type(3'b001);	// Register model should be updated in reverse order.

		    end //}

	KEEP_ALIVE : begin //{

		      lh_trans.force_drvr_oe[lane_num] = 1;

		      if (lh_trans.retrain)
		        current_cw_train_state = RETRAINING_0;
		      else if (!lh_trans.keep_alive[lane_num] & !lh_trans.retrain)
		        current_cw_train_state = TRAINED;

		      if (~bfm_or_mon)
		        update_ls1_idle3_training_type(3'b001);

		     end //}

	RETRAINING_0 : 	begin //{

		      	  lh_trans.force_drvr_oe[lane_num] = 1;

		 	  if (lh_trans.retrain_timer_done)
	         	    current_cw_train_state = RETRAIN_FAIL;
		 	  else if (!lh_trans.retrain_timer_done & !lh_trans.lane_retraining[lane_num])
	         	    current_cw_train_state = RETRAINING_1;

		      	  if (~bfm_or_mon)
		      	    update_ls1_idle3_training_type(3'b110);

	       		end //}

	RETRAINING_1 : 	begin //{

		   	  //$display($time, " : Entered SYNC_1 in lane_num %0d", lane_num);

      		      	  lh_trans.retrain_fail[lane_num] = 0;
	           	  lh_trans.retrain_lane[lane_num] = 1;

		 	  if (lh_trans.retrain_timer_done)
	         	    current_cw_train_state = RETRAIN_FAIL;
		 	  else if (!lh_trans.retrain_timer_done & lh_trans.lane_retraining[lane_num])
	         	    current_cw_train_state = RETRAINING_2;

		      	  if (~bfm_or_mon)
		      	    update_ls1_idle3_training_type(3'b110);

	       	 	end //}

	RETRAINING_2 : 	begin //{

		   	  //$display($time, " : Entered SYNC_2 in lane_num %0d", lane_num);

		 	  if (lh_trans.lane_ready[lane_num] & !lh_trans.lane_degraded[lane_num] & lh_trans.from_sc_lane_ready[lane_num])
	         	    current_cw_train_state = TRAINED;
		 	  else if ((lh_trans.retrain_timer_done & !lh_trans.retrain_timer_en) & (!lh_trans.lane_ready[lane_num] | 
					lh_trans.lane_degraded[lane_num] | !lh_trans.from_sc_lane_ready[lane_num]))
	         	    current_cw_train_state = RETRAIN_FAIL;

		      	  if (~bfm_or_mon)
		      	  begin //{
		      	    update_ls1_idle3_training_type(3'b110);
			    //if (current_cw_train_state == TRAINED)
			    //  update_ls1_idle3_cw_retraining_completed();
		      	  end //}

	       	 	end //}

	RETRAIN_FAIL : 	begin //{

      		      	  lh_trans.retrain_fail[lane_num] = 1;
      		      	  lh_trans.retrain_lane[lane_num] = 0;
      		      	  lh_trans.force_drvr_oe[lane_num] = 0;
      		      	  lh_trans.lane_trained[lane_num] = 0;

		      	  if (~bfm_or_mon)
		      	  begin //{
		      	    update_ls1_idle3_training_type(3'b110);
      		      	    update_ls1_idle3_cw_retraining_state();
		      	  end //}

		    	end //}

      endcase

      if ((prev_cw_train_state != current_cw_train_state && (current_cw_train_state == TRAINED || prev_cw_train_state == TRAINED)) && current_cw_train_state != KEEP_ALIVE && prev_cw_train_state != KEEP_ALIVE)
        `uvm_info("SRIO_LANE_HANDLER : GEN3_CW_TRAIN_SM", $sformatf(" lane_trained[%0d] is %0d Next cw train state is %0s", lane_num, lh_trans.lane_trained[lane_num], current_cw_train_state.name()), UVM_LOW)

      if (~bfm_or_mon && prev_cw_train_state != current_cw_train_state)
	current_cw_train_state_q.push_back(current_cw_train_state);

    end //}

  end //}

endtask : gen3_cw_training_sm



////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_frame_lock_sm
/// Description : Implements the frame lock state machine as defined in the 802.3-2008 specification.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_frame_lock_sm();

  bit prev_lane_trained[int];

#1;
  if (~srio_if.srio_rst_n)
  begin //{
    current_frame_lock_state = OUT_OF_FRAME;
    // questasim and vcs doesn't work properly on associatuve array methods
    // Hence, a work-around is done here by setting the array values to 1 and
    // then clearing it immediately.
    lh_trans.frame_lock[lane_num] = 1;
    lh_trans.frame_lock[lane_num] = 0;

    if (~bfm_or_mon)
      current_frame_lock_state_q.push_back(current_frame_lock_state);

  end //}

  forever
  begin //{

    prev_lane_trained[lane_num] = lh_trans.lane_trained[lane_num];

    @(negedge dme_frame_divide_clk or negedge srio_if.srio_rst_n or negedge lh_trans.lane_trained[lane_num]);

    if (~srio_if.srio_rst_n || (prev_lane_trained[lane_num] && ~lh_trans.lane_trained[lane_num]))
    begin //{

      prev_frame_lock_state = current_frame_lock_state;

      current_frame_lock_state = OUT_OF_FRAME;
      lh_trans.frame_lock[lane_num] = 0;
      new_marker = 0;

      if (~bfm_or_mon && prev_frame_lock_state != current_frame_lock_state)
        current_frame_lock_state_q.push_back(current_frame_lock_state);

    end //}
    else
    begin //{

      //`uvm_info("SRIO_LANE_HANDLER : GEN3_CW_TRAIN_SM", $sformatf(" lane_trained[%0d] is %0d Present cw train state is %0s", lane_num, lh_trans.lane_trained[lane_num], current_frame_lock_state.name()), UVM_LOW)

      prev_frame_lock_state = current_frame_lock_state;

      case (current_frame_lock_state)

	OUT_OF_FRAME : 	begin //{

      		          lh_trans.frame_lock[lane_num] = 0;
      		          new_marker = 0;

      		          current_frame_lock_state = RESET_COUNT;

		    	end //}

	RESET_COUNT : begin //{

		      	  good_markers = 0;
		      	  bad_markers = 0;

			  if (slip_done)
	      		    dme_frame_s2p_lock = 0;

		      	  slip_done = 0;

		      	  current_frame_lock_state = GET_NEW_MARKER;

		      end //}

	GET_NEW_MARKER : begin //{

		      	  frame_offset = 0;

		      	  if (new_marker)
		      	    current_frame_lock_state = TEST_MARKER;

		    	 end //}

	TEST_MARKER : begin //{

      		      	new_marker = 0;

			if (frame_marker_data == 32'hFFFF_0000) // Implies marker_valid is '1'.
			begin //{
      		      	  good_markers++;
      		      	  bad_markers = 0;
		      	  current_frame_lock_state = VALID_MARKER;
			end //}
			else
			begin //{
		      	  bad_markers++;
		      	  good_markers = 0;
		      	  current_frame_lock_state = INVALID_MARKER;
			end //}

		      end //}

	VALID_MARKER : begin //{

		      	 if ((good_markers < 2) & frame_offset)
		      	   current_frame_lock_state = GET_NEW_MARKER;
		      	 else if (good_markers == 2)
		      	   current_frame_lock_state = IN_FRAME;

		       end //}

	IN_FRAME : begin //{

		      lh_trans.frame_lock[lane_num] = 1;

		      if (frame_offset)
		        current_frame_lock_state = RESET_COUNT;

		   end //}

	INVALID_MARKER : begin //{

		 	  if ((bad_markers == 5) | (!lh_trans.frame_lock[lane_num]))
	         	    current_frame_lock_state = SLIP;
		 	  else if ((bad_markers < 5) & lh_trans.frame_lock[lane_num] & frame_offset)
	         	    current_frame_lock_state = GET_NEW_MARKER;

	       		 end //}

	SLIP : begin //{

      		 lh_trans.frame_lock[lane_num] = 0;
                 parallel_slide_mode=0;
                 note_bit_2=66;

		 if (slip_done)
	           current_frame_lock_state = RESET_COUNT;

	       end //}

      endcase

      //if (prev_frame_lock_state != current_frame_lock_state && (current_frame_lock_state == IN_FRAME || prev_frame_lock_state == IN_FRAME))
      //  `uvm_info("SRIO_LANE_HANDLER : GEN3_CW_TRAIN_SM", $sformatf(" frame_lock[%0d] is %0d Next frame lock state is %0s", lane_num, lh_trans.frame_lock[lane_num], current_frame_lock_state.name()), UVM_LOW)
      if (~bfm_or_mon && prev_frame_lock_state != current_frame_lock_state)
        current_frame_lock_state_q.push_back(current_frame_lock_state);

    end //}

  end //}

endtask : gen3_frame_lock_sm





////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : dme_wait_timer_method
/// Description : When dme_wait_timer_en is set in ~mon_type, it counts the no. of frames being
/// received by this monitor, and sets the dme_wait_timer_done for ~mon_type.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::dme_wait_timer_method();

  int local_frame_count;

  lh_common_mon_trans.dme_wait_timer_en[~mon_type][lane_num] = 1;
  lh_common_mon_trans.dme_wait_timer_en[~mon_type][lane_num] = 0;

  lh_common_mon_trans.dme_wait_timer_done[~mon_type][lane_num] = 1;
  lh_common_mon_trans.dme_wait_timer_done[~mon_type][lane_num] = 0;

  forever begin //{

    wait (lh_common_mon_trans.dme_wait_timer_en[~mon_type][lane_num] == 1);

    while (local_frame_count != lh_config.dme_wait_timer_frame_cnt)
    begin //{

      wait (frame_offset_achieved == 1);

      local_frame_count++;

      wait (frame_offset_achieved == 0);

    end //}

    local_frame_count = 0;
    lh_common_mon_trans.dme_wait_timer_done[~mon_type][lane_num] = 1;

    wait (lh_common_mon_trans.dme_wait_timer_en[~mon_type][lane_num] == 0);

    lh_common_mon_trans.dme_wait_timer_done[~mon_type][lane_num] = 0;

  end //}

endtask : dme_wait_timer_method







////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : gen3_dme_training_sm
/// Description : Implements the DME training / long-run training state machine as defined in the 
/// GEN3.0 specification.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::gen3_dme_training_sm();

#1;
  if (~srio_if.srio_rst_n)
  begin //{
    current_dme_train_state = UNTRAINED;
    // questasim and vcs doesn't work properly on associatuve array methods
    // Hence, a work-around is done here by setting the array values to 1 and
    // then clearing it immediately.
    lh_trans.lane_trained[lane_num] = 1;
    lh_trans.lane_trained[lane_num] = 0;

    lh_trans.dme_wait_timer_en[lane_num] = 1;
    lh_trans.dme_wait_timer_en[lane_num] = 0;

    lh_trans.dme_wait_timer_done[lane_num] = 1;
    lh_trans.dme_wait_timer_done[lane_num] = 0;

    lh_trans.from_dme_rcvr_ready[lane_num] = 1;
    //lh_trans.from_dme_rcvr_ready[lane_num] = 0; // Temp comment. Need to uncomment when dme training support is added in tx path

    lh_trans.current_dme_train_state[lane_num] = current_dme_train_state;

    if (~bfm_or_mon)
      current_dme_train_state_q.push_back(current_dme_train_state);

  end //}

  forever
  begin //{

    if (current_dme_train_state == CW_TRAINING_0 || current_dme_train_state == TRAINED)
    begin //{
      // just a small delay added here, so that current_cw_train_state changes from UNTRAINED state to current_dme_train_state.
      repeat(2) @(negedge dme_frame_divide_clk);
      lh_trans.dme_mode[lane_num]=0;
      wait(current_cw_train_state == UNTRAINED);
      current_dme_train_state = current_cw_train_state;

      if (~bfm_or_mon)
        update_ls1_idle3_training_type(3'b000);

      lh_trans.current_dme_train_state[lane_num] = current_dme_train_state;

      if (~bfm_or_mon)
        current_dme_train_state_q.push_back(current_dme_train_state);

    end //}

    wait (lh_trans.frame_lock[lane_num] == 1 || lh_trans.cw_lock[lane_num] == 1);

    // Since dme_frame_divide_clk will not be generated when link partner is not transmitting
    // frames. So, added divide_clk in the below sensitivity list.
    if (lh_trans.frame_lock[lane_num] == 1)
      @(negedge dme_frame_divide_clk or negedge srio_if.srio_rst_n);
    else if (lh_trans.cw_lock[lane_num] == 1)
      @(negedge divide_clk or negedge srio_if.srio_rst_n);

    if (~srio_if.srio_rst_n || (lh_trans.current_init_state == SILENT))
    begin //{

      prev_dme_train_state = current_dme_train_state;

      current_dme_train_state = UNTRAINED;
      lh_trans.force_drvr_oe[lane_num] = 0;
      lh_trans.dme_mode[lane_num] = 1;
      lh_trans.train_lane[lane_num] = 0;
      lh_trans.retrain_lane[lane_num] = 0;
      lh_trans.train_timer_en[lane_num] = 0;

      lh_trans.lane_trained[lane_num] = 0;

      lh_trans.current_dme_train_state[lane_num] = current_dme_train_state;

      if (~bfm_or_mon && prev_dme_train_state != current_dme_train_state)
        current_dme_train_state_q.push_back(current_dme_train_state);

      if (~bfm_or_mon)
        update_ls1_idle3_training_type(3'b000);

    end //}
    else
    begin //{

      //`uvm_info("SRIO_LANE_HANDLER : GEN3_CW_TRAIN_SM", $sformatf(" lane_trained[%0d] is %0d Present cw train state is %0s", lane_num, lh_trans.lane_trained[lane_num], current_dme_train_state.name()), UVM_LOW)

      prev_dme_train_state = current_dme_train_state;

      case (current_dme_train_state)

	UNTRAINED : begin //{

      		      lh_trans.force_drvr_oe[lane_num] = 0;
      		      lh_trans.dme_mode[lane_num] = 1;
      		      lh_trans.train_lane[lane_num] = 0;
      		      lh_trans.retrain_lane[lane_num] = 0;
      		      lh_trans.train_timer_en[lane_num] = 0;

		      lh_trans.xmt_equalizer = "LR_initialize";

		      if (lh_trans.drvr_oe[lane_num] & lh_trans.lane_sync[lane_num] & !lh_trans.frame_lock[lane_num])
		      begin //{
      			current_dme_train_state = CW_TRAINING_0;
		      end //}
		      else if (lh_trans.drvr_oe[lane_num] & !lh_trans.lane_sync[lane_num] & lh_trans.frame_lock[lane_num])
		      begin //{
      			current_dme_train_state = DME_TRAINING_0;
		      end //}

      		      if (~bfm_or_mon)
      		        update_ls1_idle3_training_type(3'b000);

		    end //}

	DME_TRAINING_0 : begin //{

		      	  lh_trans.train_timer_en[lane_num] = 1;

		      	  if (lh_trans.train_timer_done[lane_num])
		      	    current_dme_train_state = DME_TRAINING_FAIL;
		      	  else if (!lh_trans.train_timer_done[lane_num] & !lh_trans.lane_trained[lane_num])
		      	    current_dme_train_state = DME_TRAINING_1;

      		      	  if (~bfm_or_mon)
      		      	    update_ls1_idle3_training_type(3'b100);

		    	 end //}

	DME_TRAINING_1 : begin //{

      		      	  lh_trans.training_fail[lane_num] = 0;
		      	  lh_trans.train_lane[lane_num] = 1;

		      	  if (lh_trans.train_timer_done[lane_num])
		      	    current_dme_train_state = DME_TRAINING_FAIL;
		      	  else if (!lh_trans.train_timer_done[lane_num] & !lh_trans.drvr_oe[lane_num])
		      	    current_dme_train_state = UNTRAINED;
		      	  else if (!lh_trans.train_timer_done[lane_num] & lh_trans.drvr_oe[lane_num] & lh_trans.frame_lock[lane_num]
					& lh_trans.lane_trained[lane_num] & lh_trans.from_dme_rcvr_ready[lane_num])
		      	    current_dme_train_state = DME_TRAINING_2;

      		      	  if (~bfm_or_mon)
      		      	    update_ls1_idle3_training_type(3'b100);

		    	 end //}

	DME_TRAINING_2 : begin //{

			  if (bfm_or_mon)
      		      	    lh_trans.dme_wait_timer_en[lane_num] = 1;
			  else
			    lh_common_mon_trans.dme_wait_timer_en[mon_type][lane_num] = 1;

		      	  if (bfm_or_mon && lh_trans.dme_wait_timer_done[lane_num] & lh_trans.from_dme_rcvr_ready[lane_num])
		      	    current_dme_train_state = TRAINED;
		      	  else if (~bfm_or_mon && lh_common_mon_trans.dme_wait_timer_done[mon_type][lane_num] & lh_trans.from_dme_rcvr_ready[lane_num])
		      	    current_dme_train_state = TRAINED;
		      	  else if (!lh_trans.from_dme_rcvr_ready[lane_num])
		      	    current_dme_train_state = DME_TRAINING_1;

      		      	  if (~bfm_or_mon)
			  begin //{
      		      	    update_ls1_idle3_training_type(3'b100);
			    //if (current_dme_train_state == TRAINED)
      		      	    //   update_ls1_idle3_dme_training_completed();
			  end //}

		    	 end //}

	DME_TRAINING_FAIL : begin //{

      		      	     lh_trans.training_fail[lane_num] = 1;
		      	     current_dme_train_state = UNTRAINED;

      		      	     if (~bfm_or_mon)
			     begin //{
      		      	       update_ls1_idle3_training_type(3'b100);
      		      	       update_ls1_idle3_dme_training_state();
			     end //}

		           end //}

      endcase

      lh_trans.current_dme_train_state[lane_num] = current_dme_train_state;

      if (prev_dme_train_state != current_dme_train_state && (current_dme_train_state == TRAINED || prev_dme_train_state == TRAINED))
        `uvm_info("SRIO_LANE_HANDLER : GEN3_DME_TRAIN_SM", $sformatf(" lane_trained[%0d] is %0d Next dme train state is %0s", lane_num, lh_trans.lane_trained[lane_num], current_dme_train_state.name()), UVM_LOW)

      if (~bfm_or_mon && prev_dme_train_state != current_dme_train_state)
        current_dme_train_state_q.push_back(current_dme_train_state);

    end //}

  end //}

endtask : gen3_dme_training_sm




task srio_pl_lane_handler::comma_char_freq_check();

  int char_cnt_for_k;
  int exp_clk_comp_rate;

  if (~bfm_or_mon && ~report_error)
    exp_clk_comp_rate = lh_config.clk_compensation_seq_rate;
  if (~bfm_or_mon && report_error)
    exp_clk_comp_rate = 5000;

  forever begin //{

    @(negedge divide_clk or negedge s2p_lock);

    if (~s2p_lock)
      char_cnt_for_k = 0;

    wait(s2p_lock == 1);

    if (lh_env_config.srio_mode != SRIO_GEN30)
    begin //{

      if (lane_data_ins.character != SRIO_K || !lane_data_ins.cntl)
      begin //{
        char_cnt_for_k++;
      end //}
      else
      begin //{
        char_cnt_for_k = 0;
      end //}

      if (char_cnt_for_k > exp_clk_comp_rate)
      begin //{
        `uvm_error("SRIO_PL_LANE_HANDLER : CG_BETWEEN_CLK_COMP_CHECK", $sformatf(" Spec reference 4.7.1. Lane number : %0d. Number of code groups without a clock compensation sequences exceeded the exected count of %0d", lane_num, exp_clk_comp_rate))
        char_cnt_for_k = 0;
      end //}

    end //}
    else if (lh_env_config.srio_mode == SRIO_GEN30)
    begin //{

      if (lane_data_ins.brc3_cntl_cw_type != SKIP_MARKER)
      begin //{
        char_cnt_for_k++;
      end //}
      else
      begin //{
        char_cnt_for_k = 0;
      end //}

      if (char_cnt_for_k > exp_clk_comp_rate)
      begin //{
        `uvm_error("SRIO_PL_LANE_HANDLER : CG_BETWEEN_SKIP_MARKER_CHECK", $sformatf(" Spec reference 4.7.1. Lane number : %0d. Number of code words without a skip marker control codeword exceeded the exected count of %0d", lane_num, exp_clk_comp_rate))
        char_cnt_for_k = 0;
      end //}

    end //}
    
  end //}

endtask : comma_char_freq_check





////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : lc_cw_bip_calc_method
/// Description : This method calculates the BIP23 value of each codeword received, and also checks
/// the value against the BIP23 value of received lane check control codeword. The BIP23 value is
/// reset whenever codeword lock is lost and it is reloaded with the first lane check control
/// codeword received after codeword lock is acheived. 
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::lc_cw_bip_calc_method();
  if (~lh_trans.cw_lock[lane_num])
  begin //{
    bip23_value = 23'h00_0000;
    lc_after_cw_lock_detected = 0;
  end //}
  else if (lh_trans.cw_lock[lane_num] && ~lc_after_cw_lock_detected)
  begin //{
    if (lane_data_ins.brc3_cntl_cw_type == LANE_CHECK)
    begin //{
      bip23_value = lane_data_ins.brc3_cw[0:22];
      if(lane_data_ins.brc3_cw[0:22]==!lane_data_ins.brc3_cw[41:63])
       begin//{
        lc_after_cw_lock_detected = 1;
        `uvm_info("SRIO_LANE_HANDLER :",$sformatf("First Correct Lane Check Codeword Detected"),UVM_LOW)
        lane_data_ins.brc3_cg[3:25]=0;
        temp_bip23_value[0] = lane_data_ins.brc3_cg[21] ^ lane_data_ins.brc3_cg[44];
        for (int bip_calc=1; bip_calc<22; bip_calc++)
        begin //{
          temp_bip23_value[bip_calc] = lane_data_ins.brc3_cg[bip_calc-1] ^ lane_data_ins.brc3_cg[bip_calc+21] ^ lane_data_ins.brc3_cg[bip_calc+44];
        end //}
        temp_bip23_value[22] = lane_data_ins.brc3_cg[43] ^ lane_data_ins.brc3_cg[66];
        bip23_value = temp_bip23_value ^ bip23_value;
       end //}
    end//}

  end //}
  else if (lc_after_cw_lock_detected)
  begin //{
    if (lane_data_ins.brc3_cntl_cw_type != LANE_CHECK && lane_data_ins.brc3_cntl_cw_type != SKIP_MARKER && lane_data_ins.brc3_cntl_cw_type != SKIP)
    begin //{
      temp_bip23_value[0] = lane_data_ins.brc3_cg[21] ^ lane_data_ins.brc3_cg[44];
      for (int bip_calc=1; bip_calc<22; bip_calc++)
      begin //{
	temp_bip23_value[bip_calc] = lane_data_ins.brc3_cg[bip_calc-1] ^ lane_data_ins.brc3_cg[bip_calc+21] ^ lane_data_ins.brc3_cg[bip_calc+44];
      end //}
      temp_bip23_value[22] = lane_data_ins.brc3_cg[43] ^ lane_data_ins.brc3_cg[66];
      bip23_value = temp_bip23_value ^ bip23_value;
    end //}
    else if (lane_data_ins.brc3_cntl_cw_type == LANE_CHECK)
    begin //{
      if (lane_data_ins.brc3_cw[0:22] != bip23_value)	
      begin //{
	-> lh_trans.lanechk_cw_corrupt_bip;
        `uvm_error("SRIO_PL_LANE_HANDLER : LANE_CHECK_CW_BIP23_VALUE_CHECK", $sformatf(" Spec reference 5.5.3.2. Lane number : %0d. Incorrect BIP23 value in the received lane check control codeword. Received value is %0h, Expected value is %0h", lane_num, lane_data_ins.brc3_cw[0:22], bip23_value))
      end //}
      else
      begin //{
	-> lh_trans.lanechk_cw_correct_bip;
      end //}
      if (lane_data_ins.brc3_cw[41:63] != ~bip23_value)	
      begin //{
	-> lh_trans.lanechk_cw_corrupt_bip;
        `uvm_error("SRIO_PL_LANE_HANDLER : LANE_CHECK_CW_iBIP23_VALUE_CHECK", $sformatf(" Spec reference 5.5.3.2. Lane number : %0d. Incorrect iBIP23 value in the received lane check control codeword. Received value is %0h, Expected value is %0h", lane_num, lane_data_ins.brc3_cw[41:63], ~bip23_value))
      end //}
      if ({lane_data_ins.brc3_cw[23:29], lane_data_ins.brc3_cw[36:40]} != 12'hB55)	
      begin //{
	-> lh_trans.lanechk_cw_corrupt_bip;
        `uvm_error("SRIO_PL_LANE_HANDLER : LANE_CHECK_CW_FIXED_VALUE_CHECK", $sformatf(" Spec reference 5.5.3.2. Lane number : %0d. Incorrect fixed value in the received lane check control codeword. Received value is %0h, Expected value is 12'hB55", lane_num, {lane_data_ins.brc3_cw[23:29], lane_data_ins.brc3_cw[36:40]}))
      end //}
      bip23_value = lane_data_ins.brc3_cw[0:22];
      bip23_value = 0; 
      temp_bip23_value=0;
      lane_data_ins.brc3_cg[3:25]=0;
      temp_bip23_value[0] = lane_data_ins.brc3_cg[21] ^ lane_data_ins.brc3_cg[44];
      for (int bip_calc=1; bip_calc<22; bip_calc++)
      begin //{
        temp_bip23_value[bip_calc] = lane_data_ins.brc3_cg[bip_calc-1] ^ lane_data_ins.brc3_cg[bip_calc+21] ^ lane_data_ins.brc3_cg[bip_calc+44];
      end //}
      temp_bip23_value[22] = lane_data_ins.brc3_cg[43] ^ lane_data_ins.brc3_cg[66];
      bip23_value = temp_bip23_value ^ bip23_value;
    end //}
  end //}
endtask : lc_cw_bip_calc_method
////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_ls1_idle3_training_type
/// Description : This method updates the IDLE3 Training Type field of LaneN_Status_1 CSR.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_ls1_idle3_training_type(bit [2:0] training_type_val);

  if (lane_num == 0)
    void'(lh_reg_model.Lane_0_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 1)
    void'(lh_reg_model.Lane_1_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 2)
    void'(lh_reg_model.Lane_2_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 3)
    void'(lh_reg_model.Lane_3_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 4)
    void'(lh_reg_model.Lane_4_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 5)
    void'(lh_reg_model.Lane_5_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 6)
    void'(lh_reg_model.Lane_6_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 7)
    void'(lh_reg_model.Lane_7_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 8)
    void'(lh_reg_model.Lane_8_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 9)
    void'(lh_reg_model.Lane_9_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 10)
    void'(lh_reg_model.Lane_10_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 11)
    void'(lh_reg_model.Lane_11_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 12)
    void'(lh_reg_model.Lane_12_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 13)
    void'(lh_reg_model.Lane_13_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 14)
    void'(lh_reg_model.Lane_14_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));
  else if (lane_num == 15)
    void'(lh_reg_model.Lane_15_Status_1_CSR.IDLE3_Training_Type.predict(training_type_val));

endtask : update_ls1_idle3_training_type




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_ls1_idle3_dme_training_state
/// Description : This method updates the IDLE3 DME Training state field of LaneN_Status_1 CSR.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_ls1_idle3_dme_training_state();

  if (lane_num == 0)
    void'(lh_reg_model.Lane_0_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 1)
    void'(lh_reg_model.Lane_1_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 2)
    void'(lh_reg_model.Lane_2_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 3)
    void'(lh_reg_model.Lane_3_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 4)
    void'(lh_reg_model.Lane_4_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 5)
    void'(lh_reg_model.Lane_5_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 6)
    void'(lh_reg_model.Lane_6_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 7)
    void'(lh_reg_model.Lane_7_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 8)
    void'(lh_reg_model.Lane_8_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 9)
    void'(lh_reg_model.Lane_9_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 10)
    void'(lh_reg_model.Lane_10_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 11)
    void'(lh_reg_model.Lane_11_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 12)
    void'(lh_reg_model.Lane_12_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 13)
    void'(lh_reg_model.Lane_13_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 14)
    void'(lh_reg_model.Lane_14_Status_1_CSR.IDLE3_DME_Training_State.predict(1));
  else if (lane_num == 15)
    void'(lh_reg_model.Lane_15_Status_1_CSR.IDLE3_DME_Training_State.predict(1));

endtask : update_ls1_idle3_dme_training_state




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_ls1_idle3_cw_training_state
/// Description : This method updates the IDLE3 SC Training state field of LaneN_Status_1 CSR.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_ls1_idle3_cw_training_state();

  if (lane_num == 0)
    void'(lh_reg_model.Lane_0_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 1)
    void'(lh_reg_model.Lane_1_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 2)
    void'(lh_reg_model.Lane_2_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 3)
    void'(lh_reg_model.Lane_3_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 4)
    void'(lh_reg_model.Lane_4_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 5)
    void'(lh_reg_model.Lane_5_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 6)
    void'(lh_reg_model.Lane_6_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 7)
    void'(lh_reg_model.Lane_7_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 8)
    void'(lh_reg_model.Lane_8_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 9)
    void'(lh_reg_model.Lane_9_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 10)
    void'(lh_reg_model.Lane_10_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 11)
    void'(lh_reg_model.Lane_11_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 12)
    void'(lh_reg_model.Lane_12_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 13)
    void'(lh_reg_model.Lane_13_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 14)
    void'(lh_reg_model.Lane_14_Status_1_CSR.IDLE3_SC_Training_State.predict(1));
  else if (lane_num == 15)
    void'(lh_reg_model.Lane_15_Status_1_CSR.IDLE3_SC_Training_State.predict(1));

endtask : update_ls1_idle3_cw_training_state




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_ls1_idle3_cw_retraining_state
/// Description : This method updates the IDLE3 SC Re-Training state field of LaneN_Status_1 CSR.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_ls1_idle3_cw_retraining_state();

  if (lane_num == 0)
    void'(lh_reg_model.Lane_0_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 1)
    void'(lh_reg_model.Lane_1_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 2)
    void'(lh_reg_model.Lane_2_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 3)
    void'(lh_reg_model.Lane_3_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 4)
    void'(lh_reg_model.Lane_4_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 5)
    void'(lh_reg_model.Lane_5_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 6)
    void'(lh_reg_model.Lane_6_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 7)
    void'(lh_reg_model.Lane_7_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 8)
    void'(lh_reg_model.Lane_8_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 9)
    void'(lh_reg_model.Lane_9_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 10)
    void'(lh_reg_model.Lane_10_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 11)
    void'(lh_reg_model.Lane_11_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 12)
    void'(lh_reg_model.Lane_12_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 13)
    void'(lh_reg_model.Lane_13_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 14)
    void'(lh_reg_model.Lane_14_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));
  else if (lane_num == 15)
    void'(lh_reg_model.Lane_15_Status_1_CSR.IDLE3_SC_Retraining_State.predict(1));

endtask : update_ls1_idle3_cw_retraining_state




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_ls2_reg
/// Description : This method updates the Lane N Status 2 CSR.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_ls2_reg();

  if (lane_num == 0)
    void'(lh_reg_model.Lane_0_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 1)
    void'(lh_reg_model.Lane_1_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 2)
    void'(lh_reg_model.Lane_2_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 3)
    void'(lh_reg_model.Lane_3_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 4)
    void'(lh_reg_model.Lane_4_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 5)
    void'(lh_reg_model.Lane_5_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 6)
    void'(lh_reg_model.Lane_6_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 7)
    void'(lh_reg_model.Lane_7_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 8)
    void'(lh_reg_model.Lane_8_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 9)
    void'(lh_reg_model.Lane_9_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 10)
    void'(lh_reg_model.Lane_10_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 11)
    void'(lh_reg_model.Lane_11_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 12)
    void'(lh_reg_model.Lane_12_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 13)
    void'(lh_reg_model.Lane_13_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 14)
    void'(lh_reg_model.Lane_14_Status_2_CSR.predict(ls2_reg_val));
  else if (lane_num == 15)
    void'(lh_reg_model.Lane_15_Status_2_CSR.predict(ls2_reg_val));

endtask : update_ls2_reg




////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_ls3_reg
/// Description : This method updates the Lane N Status 3 CSR.
////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_ls3_reg();

  if (lane_num == 0)
    void'(lh_reg_model.Lane_0_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 1)
    void'(lh_reg_model.Lane_1_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 2)
    void'(lh_reg_model.Lane_2_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 3)
    void'(lh_reg_model.Lane_3_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 4)
    void'(lh_reg_model.Lane_4_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 5)
    void'(lh_reg_model.Lane_5_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 6)
    void'(lh_reg_model.Lane_6_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 7)
    void'(lh_reg_model.Lane_7_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 8)
    void'(lh_reg_model.Lane_8_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 9)
    void'(lh_reg_model.Lane_9_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 10)
    void'(lh_reg_model.Lane_10_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 11)
    void'(lh_reg_model.Lane_11_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 12)
    void'(lh_reg_model.Lane_12_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 13)
    void'(lh_reg_model.Lane_13_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 14)
    void'(lh_reg_model.Lane_14_Status_3_CSR.predict(ls3_reg_val));
  else if (lane_num == 15)
    void'(lh_reg_model.Lane_15_Status_3_CSR.predict(ls3_reg_val));

endtask : update_ls3_reg




//////////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name : update_error_detect_csr
/// Description : This method updates the Port n Error detect CSR when lane specific errors are detected.
/// It also checks if corresponding bit is set in error rate CSR, and updates the error rate counter in 
/// Error Rate CSR.
//////////////////////////////////////////////////////////////////////////////////////////////////////////
task srio_pl_lane_handler::update_error_detect_csr(string csr_field_name);

  bit error_enable;
  bit [7:0] error_rate_counter;

  if (csr_field_name == "INVALID_CHAR")
  begin //{
    register_update_method("Error_Detect_CSR", "Received_illegal_or_invalid_character", 64, "lh_reg_model", reqd_field_name["Received_illegal_or_invalid_character"]);
    void'(reqd_field_name["Received_illegal_or_invalid_character"].predict(1));
    //void'(lh_reg_model.Port_0_Error_Detect_CSR.Received_illegal_or_invalid_character.predict(1));
    register_update_method("Error_Rate_Enable_CSR", "Received_illegal_or_invalid_character_enable", 64, "lh_reg_model", reqd_field_name["Received_illegal_or_invalid_character_enable"]);
    error_enable = reqd_field_name["Received_illegal_or_invalid_character_enable"].get();
    //error_enable = lh_reg_model.Port_0_Error_Rate_Enable_CSR.Received_illegal_or_invalid_character_enable.get();
    register_update_method("Error_Detect_CSR", "Delineation_error", 64, "lh_reg_model", reqd_field_name["Delineation_error"]);
    void'(reqd_field_name["Delineation_error"].predict(1));
    //void'(lh_reg_model.Port_0_Error_Detect_CSR.Delineation_error.predict(1));	// Delin error will be set when invalid_cg is detected.
    if (~error_enable)
    begin //{
      register_update_method("Error_Rate_Enable_CSR", "Delineation_error_enable", 64, "lh_reg_model", reqd_field_name["Delineation_error_enable"]);
      error_enable = reqd_field_name["Delineation_error_enable"].get();
      //error_enable = lh_reg_model.Port_0_Error_Rate_Enable_CSR.Delineation_error_enable.get();	// Checking error_enable only if it is not set before.
    end //}
  end //}
  else if (csr_field_name == "DESCR_SYNC_LOSS")
  begin //{
    register_update_method("Error_Detect_CSR", "Loss_of_descrambler_synchronization", 64, "lh_reg_model", reqd_field_name["Loss_of_descrambler_synchronization"]);
    void'(reqd_field_name["Loss_of_descrambler_synchronization"].predict(1));
    //void'(lh_reg_model.Port_0_Error_Detect_CSR.Loss_of_descrambler_synchronization.predict(1));
    register_update_method("Error_Rate_Enable_CSR", "Loss_of_descrambler_synchronization_enable", 64, "lh_reg_model", reqd_field_name["Loss_of_descrambler_synchronization_enable"]);
    error_enable = reqd_field_name["Loss_of_descrambler_synchronization_enable"].get();
    //error_enable = lh_reg_model.Port_0_Error_Rate_Enable_CSR.Loss_of_descrambler_synchronization_enable.get();
  end //}
  else if (csr_field_name == "DELIN_ERR")
  begin //{
    register_update_method("Error_Detect_CSR", "Delineation_error", 64, "lh_reg_model", reqd_field_name["Delineation_error"]);
    void'(reqd_field_name["Delineation_error"].predict(1));
    //void'(lh_reg_model.Port_0_Error_Detect_CSR.Delineation_error.predict(1));
    register_update_method("Error_Rate_Enable_CSR", "Delineation_error_enable", 64, "lh_reg_model", reqd_field_name["Delineation_error_enable"]);
    error_enable = reqd_field_name["Delineation_error_enable"].get();
    //error_enable = lh_reg_model.Port_0_Error_Rate_Enable_CSR.Delineation_error_enable.get();
  end //}
  //else if (csr_field_name == "INVALID_OS")
  //begin //{
  //  void'(lh_reg_model.Port_0_Error_Detect_CSR.Invalid_ordered_sequence.predict(1));
  //  error_enable = lh_reg_model.Port_0_Error_Rate_Enable_CSR.Invalid_ordered_sequence_enable.get();
  //end //}

  if (error_enable)
  begin //{
    register_update_method("Error_Rate_CSR", "Error_Rate_Counter", 64, "lh_reg_model", reqd_field_name["Error_Rate_Counter"]);
    error_rate_counter = reqd_field_name["Error_Rate_Counter"].get();
    //error_rate_counter = lh_reg_model.Port_0_Error_Rate_CSR.Error_Rate_Counter.get();
    error_rate_counter = {error_rate_counter[0], error_rate_counter[1], error_rate_counter[2], error_rate_counter[3], error_rate_counter[4], error_rate_counter[5], error_rate_counter[6], error_rate_counter[7]};
    if (error_rate_counter < 8'hFF)
    begin //{
      error_rate_counter++;
      error_rate_counter = {error_rate_counter[0], error_rate_counter[1], error_rate_counter[2], error_rate_counter[3], error_rate_counter[4], error_rate_counter[5], error_rate_counter[6], error_rate_counter[7]};
      register_update_method("Error_Rate_CSR", "Error_Rate_Counter", 64, "lh_reg_model", reqd_field_name["Error_Rate_Counter"]);
      void'(reqd_field_name["Error_Rate_Counter"].predict(error_rate_counter));
      //void'(lh_reg_model.Port_0_Error_Rate_CSR.Error_Rate_Counter.predict(error_rate_counter));
    end //}
  end //}

endtask : update_error_detect_csr




////////////////////////////////////////////////////////////////////////////////////////////////////////////
/// Name :register_update_method 
/// Description : This method updates the appropriate register based on the port number configured.
/// It initially does a string concatenation based on the port number to form the register name, and then
/// gets the register name using the get_reg_by_name function. It then calculates the offset of the 
/// required register and then gets its name through get_reg_by_offset function. With the required register
/// name, the required field name is obtained from the get_field_by_name function and returned.
////////////////////////////////////////////////////////////////////////////////////////////////////////////
task automatic srio_pl_lane_handler::register_update_method(string reg_name, string field_name, int offset, string reg_ins, output uvm_reg_field out_field_name);

  string temp_reg_name;
  string reg_name_prefix;
  uvm_reg_addr_t reg_addr;
  uvm_reg reqd_reg_name;
  uvm_reg reg_name1;

  if (lh_env_config.port_number == 0)
    reg_name_prefix = "Port_0_";
  else if (lh_env_config.port_number == 1)
    reg_name_prefix = "Port_1_";
  else if (lh_env_config.port_number == 2)
    reg_name_prefix = "Port_2_";
  else if (lh_env_config.port_number == 3)
    reg_name_prefix = "Port_3_";
  else if (lh_env_config.port_number == 4)
    reg_name_prefix = "Port_4_";
  else if (lh_env_config.port_number == 5)
    reg_name_prefix = "Port_5_";
  else if (lh_env_config.port_number == 6)
    reg_name_prefix = "Port_6_";
  else if (lh_env_config.port_number == 7)
    reg_name_prefix = "Port_7_";
  else if (lh_env_config.port_number == 8)
    reg_name_prefix = "Port_8_";
  else if (lh_env_config.port_number == 9)
    reg_name_prefix = "Port_9_";
  else if (lh_env_config.port_number == 10)
    reg_name_prefix = "Port_10_";
  else if (lh_env_config.port_number == 11)
    reg_name_prefix = "Port_11_";
  else if (lh_env_config.port_number == 12)
    reg_name_prefix = "Port_12_";
  else if (lh_env_config.port_number == 13)
    reg_name_prefix = "Port_13_";
  else if (lh_env_config.port_number == 14)
    reg_name_prefix = "Port_14_";
  else if (lh_env_config.port_number == 15)
    reg_name_prefix = "Port_15_";
  else
    reg_name_prefix = "Port_0_";

  temp_reg_name = {reg_name_prefix, reg_name};

  if (reg_ins == "lh_reg_model")
    reg_name1 = lh_reg_model.get_reg_by_name(temp_reg_name);
  else if (reg_ins == "lh_reg_model_tx")
    reg_name1 = lh_env_config.srio_reg_model_tx.get_reg_by_name(temp_reg_name);
  else if (reg_ins == "lh_reg_model_rx")
    reg_name1 = lh_env_config.srio_reg_model_rx.get_reg_by_name(temp_reg_name);

  if (reg_name1 == null)
    `uvm_warning("NULL_REGISTER_ACCESS", $sformatf(" No register found with name %0s", temp_reg_name))
  reg_addr = reg_name1.get_offset();

  if (lh_env_config.srio_mode != SRIO_GEN30 && lh_env_config.spec_support != V30)
  begin //{
    if (reg_name == "Link_Maintenance_Response_CSR" || reg_name == "Control_2_CSR" || reg_name == "Error_and_Status_CSR" || reg_name == "Control_CSR")
      offset = 32;
  end //}

  if (reg_ins == "lh_reg_model")
    reqd_reg_name = lh_reg_model.srio_reg_block_map.get_reg_by_offset(reg_addr+(lh_env_config.port_number*offset));
  else if (reg_ins == "lh_reg_model_tx")
    reqd_reg_name = lh_env_config.srio_reg_model_tx.srio_reg_block_map.get_reg_by_offset(reg_addr+(lh_env_config.port_number*offset));
  else if (reg_ins == "lh_reg_model_rx")
    reqd_reg_name = lh_env_config.srio_reg_model_rx.srio_reg_block_map.get_reg_by_offset(reg_addr+(lh_env_config.port_number*offset));

  if (reqd_reg_name == null)
    `uvm_warning("NULL_REGISTER_ACCESS", $sformatf(" Register %0s. Base address : %0h, Accessed address : %0h", temp_reg_name, reg_addr, reg_addr+(lh_env_config.port_number*offset)))
  else
  begin //{
    out_field_name = reqd_reg_name.get_field_by_name(field_name);
  end //}

endtask : register_update_method
