
////////////////////////////////////////////////////////////////////////////////
//(c) Copyright 2013 Mobiveil, Inc. All rights reserved
//
// File    :  srio_ll_lfc_xon_test.sv
// Project :  srio vip
// Purpose :  LFC Test 
// Author  :  Mobiveil
//
// Test for LFC with XON Only
//
////////////////////////////////////////////////////////////////////////////////

class srio_ll_lfc_xon_test extends srio_base_test;

  `uvm_component_utils(srio_ll_lfc_xon_test)

  srio_ll_lfc_xon_seq lfc_xon_seq;
    
  function new(string name, uvm_component parent=null);
    super.new(name, parent);
  endfunction

    task run_phase( uvm_phase phase );
    super.run_phase(phase);
    lfc_xon_seq = srio_ll_lfc_xon_seq::type_id::create("lfc_xon_seq");

    phase.raise_objection( this );
    lfc_xon_seq.start( env1.e_virtual_sequencer);

    #2000ns;
       phase.drop_objection(this);
    
  endtask


endclass


