//=============================================================================
//== (c) Copyright 2013 Mobiveil Inc. All rights reserved
//== File       : srio_test_lib_pkg.sv
//== Project    : srio vip
//== Author     : Mobiveil
//== Purpose    :
//==  Package for created tests.
//==
//==
//==
//==============================================================================

package srio_test_lib_pkg;
`include "uvm_macros.svh"

import uvm_pkg::*;
import srio_env_pkg::*;
import srio_seq_lib_pkg::*;

`include "srio_pl_test_cb.sv"
`include "srio_base_test.sv"
`include "srio_ll_test_cb.sv"
`include "srio_tl_test_cb.sv"
`include "srio_ll_default_test.sv"
`include "srio_ll_nread_req_test.sv"
`include "srio_ll_message_random_test.sv"
`include "srio_ll_atomic_inc_test.sv"
`include "srio_ll_atomic_dec_test.sv"
`include "srio_ll_atomic_set_test.sv"
`include "srio_ll_atomic_clear_test.sv"
`include "srio_ll_nwrite_req_test.sv"
`include "srio_ll_nwrite_r_req_test.sv"
`include "srio_ll_atomic_swap_test.sv"
`include "srio_ll_atomic_compare_and_swap_test.sv"
`include "srio_ll_atomic_test_and_swap_test.sv"
`include "srio_ll_swrite_req_test.sv"
`include "srio_ll_maintenance_rd_req_test.sv"
`include "srio_ll_maintenance_wr_req_test.sv"
`include "srio_ll_maintenance_rd_resp_req_test.sv"
`include "srio_ll_maintenance_wr_resp_req_test.sv"
`include "srio_ll_maintenance_port_wr_req_test.sv"
`include "srio_ll_doorbell_req_test.sv"
`include "srio_ll_msg_ssize_8byte_req_test.sv"
`include "srio_ll_msg_ssize_16byte_req_test.sv"
`include "srio_ll_msg_ssize_32byte_req_test.sv"
`include "srio_ll_msg_ssize_64byte_req_test.sv"
`include "srio_ll_msg_ssize_128byte_req_test.sv"
`include "srio_ll_msg_ssize_256byte_req_test.sv"
`ifdef SRIO_VIP_B2B
`include "srio_ll_lfc_prio_lesser_ds_xon_xoff_test.sv"
`include "srio_ll_lfc_prio_ds_block_release_xon_xoff_test.sv"
`include "srio_ll_lfc_ds_random_prio_xon_xoff_test.sv"
`include "srio_ll_lfc_orphaned_xoff_test.sv"
`include "srio_ll_lfc_user_gen_xon_xoff_test.sv"
`include "srio_ll_lfc_xon_xoff_test.sv"
`include "srio_ll_lfc_multi_xon_xoff_same_flowid_test.sv"
`include "srio_ll_lfc_multi_xoff_orphaned_test.sv"
`include "srio_ll_lfc_xon_without_xoff_test.sv"
`include "srio_ll_lfc_test.sv"
`include "srio_ll_lfc_multi_xon_xoff_diff_flowid_test.sv"
`include "srio_ll_lfc_timeout_check_test.sv"
`include "srio_ll_lfc_timeout_check1_test.sv"
`include "srio_ll_lfc_random_test.sv"
`include "srio_ll_lfc_with_diff_id_test.sv"
`include "srio_ll_lfc_unsupported_flowid_test.sv"
`include "srio_ll_lfc_prio_greater_ds_xon_xoff_test.sv"
`include "srio_ll_traffic_mgmt_lfc_xoff_xon_test.sv"
`include "srio_ll_vc_ds_lfc_xoff_xon_test.sv"
`include "srio_ll_vc_support_2_lfc_xoff_xon_test.sv"
`include "srio_ll_vc_support_4_lfc_xoff_xon_test.sv"
`include "srio_ll_vc_support_8_lfc_xoff_xon_test.sv"
`include "srio_ll_vc_unsupport_flowid_ds_lfc_xoff_xon_test.sv"
`include "srio_ll_vc_support_swrite_nwrite_lfc_xoff_xon_test.sv"
`include "srio_ll_vc_support_random_ds_lfc_xoff_xon_test.sv"
`include "srio_ll_fam_req_0_spdu_xon_0_req_1_spdu_ds_spdu_xon_1_ds_spdu_test.sv"
`include "srio_ll_fam_req_0_mpdu_xon_0_ds_mpdu_xoff_0_release_0_test.sv"
`include "srio_ll_fam_req_1_mpdu_xon_1_ds_mpdu_xoff_1_release_1_test.sv"
`include "srio_ll_fam_no_req_xon_1_ds_mpdu_test.sv"
`include "srio_ll_fam_no_req_xon_0_ds_mpdu_test.sv"
`include "srio_ll_fam_no_req_xon_1_ds_spdu_test.sv"
`include "srio_ll_fam_no_req_xon_0_ds_spdu_test.sv"
`include "srio_ll_fam_no_req_no_xon_ds_mpdu_test.sv"
`include "srio_ll_fam_no_req_no_xon_ds_spdu_test.sv"
`include "srio_ll_fam_no_req_no_xon_no_ds_release_1_test.sv"
`include "srio_ll_fam_no_req_no_xon_no_ds_release_0_test.sv"
`include "srio_ll_fam_req_mpdu_no_xon_no_ds_mpdu_release_1_test.sv"
`include "srio_ll_fam_req_mpdu_no_xon_no_ds_mpdu_release_0_test.sv"
`include "srio_ll_fam_req_mpdu_xon_0_no_ds_mpdu_release_1_test.sv"
`include "srio_ll_fam_req_mpdu_xon_1_no_ds_mpdu_release_1_test.sv"
`include "srio_ll_fam_req_mpdu_xon_0_no_ds_mpdu_release_0_test.sv"
`include "srio_ll_fam_req_mpdu_xon_1_no_ds_mpdu_release_0_test.sv"
`include "srio_ll_fam_req_mpdu_xon_0_xon_0_ds_mpdu_release_0_test.sv"
`include "srio_ll_fam_req_spdu_xon_1_xon_1_ds_spdu_test.sv"
`include "srio_ll_fam_req_mpdu_xon_1_xon_1_ds_mpdu_release_1_test.sv"
`include "srio_ll_fam_req_spdu_xon_0_xon_0_ds_spdu_test.sv"
`include "srio_ll_fam_req_spdu_xon_1_xoff_1_ds_spdu_test.sv"
`include "srio_ll_fam_req_spdu_xon_0_xoff_0_ds_spdu_test.sv"
`include "srio_ll_fam_req_spdu_xon_1_ds_spdu_xoff_1_xon_1_test.sv"
`include "srio_ll_fam_req_spdu_xon_0_ds_spdu_xoff_0_xon_0_test.sv"
`include "srio_ll_fam_req_no_xon_ds_release_multi_pdu_0_test.sv"
`include "srio_ll_fam_req_no_xon_ds_release_multi_pdu_1_test.sv"
`include "srio_ll_fam_req_xoff_ds_release_multi_pdu_1_test.sv"
`include "srio_ll_fam_req_xoff_ds_release_multi_pdu_0_test.sv"
`include "srio_ll_fam_req_xon_ds_without_release_multi_pdu_1_test.sv"
`include "srio_ll_fam_req_xon_ds_without_release_multi_pdu_0_test.sv"
`include "srio_ll_fam_req_spdu_xon_ds_multi_pdu_1_test.sv"
`include "srio_ll_fam_req_spdu_xon_ds_multi_pdu_0_test.sv"
`include "srio_ll_fam_req_xon_ds_release_multi_pdu_0_test.sv"
`include "srio_ll_fam_req_xon_ds_single_pdu_0_test.sv"
`include "srio_ll_fam_req_xon_ds_release_multi_pdu_1_test.sv"
`include "srio_ll_fam_req_xon_ds_single_pdu_1_test.sv"
`include "srio_ll_fam_req_no_xon_ds_single_pdu_1_test.sv"
`include "srio_ll_fam_req_no_xon_ds_single_pdu_0_test.sv"
`include "srio_ll_fam_req_xon_ds_release_single_pdu_1_test.sv"
`include "srio_ll_fam_req_xon_ds_release_single_pdu_0_test.sv"
`include "srio_ll_fam_req_xoff_ds_single_pdu_0_test.sv"
`include "srio_ll_fam_req_xoff_ds_single_pdu_1_test.sv"
`include "srio_ll_fam_req_xon_ds_single_pdu_0_flowid_error_test.sv"
`include "srio_ll_fam_req_xon_ds_single_pdu_1_flowid_error_test.sv"
`include "srio_ll_fam_req_mpdu_xon_1_ds_mpdu_1_release_1_flowid_error_test.sv"
`include "srio_ll_fam_req_mpdu_xon_0_ds_mpdu_0_release_0_flowid_error_test.sv"
`include "srio_ll_fam_req_spdu_xon_1_ds_spdu_lesser_flowid_test.sv"
`include "srio_ll_fam_req_spdu_xon_0_ds_spdu_lesser_flowid_test.sv"
`include "srio_ll_fam_req_spdu_xon_1_ds_spdu_greater_flowid_test.sv"
`include "srio_ll_fam_req_spdu_xon_0_ds_spdu_greater_flowid_test.sv"
`include "srio_ll_fam_mpdu_xon_1_ds_mpdu_release_1_flowid_error_test.sv"
`include "srio_ll_fam_mpdu_xon_0_ds_mpdu_release_0_flowid_error_test.sv"
`include "srio_ll_fam_req_mpdu_xon_1_ds_mpdu_xoff_1_ds_mpdu_release_1_test.sv"
`include "srio_ll_fam_req_mpdu_xon_0_ds_mpdu_xoff_0_ds_mpdu_release_0_test.sv"
`include "srio_ll_ds_traffic_mgmt_basic_stream_xoff_test.sv"
`include "srio_ll_ds_traffic_mgmt_user_credit_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_user_rate_xoff_xon_test.sv"
`include "srio_ll_io_msg_gsm_ds_random_test.sv"
`include "srio_ll_ds_traffic_mgmt_user_credit_err_test.sv"
`include "srio_ll_ds_traffic_mgmt_basic_specific_stream_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_rate_specific_stream_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_credit_specific_stream_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_basic_specific_cos_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_test.sv"
`include "srio_ll_ds_traffic_mgmt_rate_specific_cos_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_credit_specific_cos_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_basic_group_of_cos_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_rate_group_of_cos_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_credit_group_of_cos_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_basic_random_cos_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_rate_random_cos_xoff_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_credit_random_cos_xoff_xon_test.sv"
`include "srio_ll_ds_all_traffic_basic_xoff_xon_test.sv"
`include "srio_ll_ds_all_traffic_rate_xoff_xon_test.sv"
`include "srio_ll_ds_all_traffic_credit_xoff_xon_test.sv"
`include "srio_pl_pkt_rty_cs_test.sv"
`include "srio_pl_pkt_na_cs_test.sv"
`include "srio_pl_asymmetry_s1xmx2_axe_test.sv"
`include "srio_pl_asymmetry_s2xmx2_axe_test.sv"
`include "srio_pl_asymmetry_s1xmx_s1xmx3_test.sv"
`include "srio_pl_asymmetry_s2xmx_s2xmx3_test.sv"
`include "srio_pl_asymmetry_xmit_width_cmd1_test.sv"
`include "srio_pl_asymmetry_rcv_width_cmd1_test.sv"
`include "srio_pl_asymmetry_sm_test.sv"
`include "srio_pl_nxm_2xm_asymmetry_sm_test.sv" 
`include "srio_pl_nxm_2xm_1xm_asymmetry_sm_test.sv"
`include "srio_pl_nxm_1xm_asymmetry_sm_test.sv"
`include "srio_pl_asymmetry_2xm_disable_1xm_test.sv" 
`include "srio_pl_asymmetry_nxm_disable_1xm_test.sv" 
`include "srio_pl_asymmetry_nxm_disable_2xm_test.sv"
`include "srio_pl_asymmetry_xmt_width_port_cmd_nx_2x_1x_nx_test.sv"
`include "srio_pl_cw_train1_untrned_test.sv"
`include "srio_pl_timestamp_check_test.sv"
`include "srio_pl_asymmetry_rcv_1x_recovery_test.sv"
`include "srio_pl_asymmetry_rcv_2x_recovery_test.sv"
`include "srio_pl_asymmetry_rcv_s2xmrcv_rwn_test.sv"
`include "srio_pl_force1x_mode_portwidth_override_test.sv"
`include "srio_pl_force1x_mode_laner_portwidth_override_test.sv"
`include "srio_pl_nxmode_enabled_2x_disabled_portwidth_override_test.sv"
`include "srio_pl_2xmode_enabled_nx_disabled_portwidth_override_test.sv"
`include "srio_pl_cw_retrain_test.sv"   
`include "srio_pl_ns1_ns2_ns_sm_test.sv"  //need to verify
`include "srio_pl_ns1_ns2_ns1_ns2_sm_test.sv" //need to verify
`include "srio_pl_pkt_flow_control_mode_transmit_test.sv"//
`include "srio_pl_diff_mode_13_21_test.sv"
`include "srio_pl_diff_mode_13_22_test.sv"
`include "srio_pl_diff_mode_22_21_test.sv"
`include "srio_ll_nread_req_env1_env2_test.sv"
`include "srio_pl_dme_min_limit_test.sv"
`include "srio_pl_dme_port_initialize_to_silent_test.sv"
`include "srio_ll_fam_pipeline_req_multi_pdu_test.sv"
`include "srio_pl_ct_mode_multi_vc_support_test.sv"  ///need to verify
`include "srio_pl_ct_mode_vc_support_transmit_mode_test.sv"
`include "srio_ll_outstanding_unack_req_test.sv"
`include "srio_ll_msg_outoforder_resp_test.sv"
`include "srio_ll_resp_error_ratio_test.sv"
`include "srio_ll_resp_no_response_ratio_test.sv"
`include "srio_ll_resp_gen_mode_test.sv"
`include "srio_ll_gsm_resp_retry_ratio_test.sv"
`include "srio_ll_msg_db_resp_retry_ratio_test.sv"
`include "srio_ll_ds_traffic_mgmt_xon_test.sv"
`include "srio_ll_ds_traffic_mgmt_tmop_err_test.sv" 
`include "srio_ll_ds_traffic_mgmt_parameter1_err_test.sv"
`include "srio_ll_ds_traffic_mgmt_xtype_err_test.sv"
`include "srio_ll_ds_traffic_mgmt_xoff_test.sv"
`include "srio_ll_msg_mseg_resp_with_payload_err_test.sv"
`include "srio_ll_msg_mseg_resp_with_invalid_status_err_test.sv"
`include "srio_ll_msg_mseg_resp_with_invalid_tgtinfo_err_test.sv"
`include "srio_ll_msg_db_resp_rand_test.sv"
`include "srio_ll_io_resp_rand_test.sv"
`include "srio_ll_gsm_resp_rand_test.sv"
`include "srio_ll_msg_mseg_resp_retry_ratio_test.sv"
`include "srio_ll_gsm_resp_err_ratio_test.sv"
`include "srio_ll_msg_resp_err_ratio_test.sv"
`include "srio_ll_msg_max_resp_delay_test.sv"
`include "srio_ll_gsm_address_collision_test.sv"
`include "srio_ll_msg_consecutive_resp_err_test.sv"
`include "srio_ll_default_illegal_resp_status_err_test.sv"
`include "srio_ll_nwrite_r_gsm_illegal_resp_err_test.sv"
`include "srio_txrx_model_test.sv"
`include "srio_pl_asymmetry_rcv_s1xmrcv_rwn_test.sv"
`include "srio_pl_cw_retrain_timeout_test.sv"
`include "srio_pl_asymmetry_rcv_s1xmrcv_are_test.sv"
`include "srio_pl_asymmetry_rcv_s2xmrcv_are_test.sv"
`include "srio_pl_asymmetry_rcv_2x_recovery_to_are_test.sv"
`include "srio_pl_asymmetry_rcv_1x_recovery_to_are_test.sv"
`include "srio_pl_force_1xmode_lane0_2x_support_test.sv"
`include "srio_pl_asymmetry_rcv_1x_mode_rcv_to_are_test.sv"
`include "srio_pl_asymmetry_rcv_2x_mode_rcv_to_are_test.sv"
`include "srio_pl_asymmetry_rcv_1xmrcv_1xmrcva_test.sv"
`include "srio_pl_asymmetry_rcv_2xmrcv_2xmrcva_test.sv"
`include "srio_pl_asymmetry_rcv_x1mrcv_x1rec_x1mrcv_test.sv"
`include "srio_pl_asymmetry_rcv_x2mrcv_x2rec_x2mrcv_test.sv"
`include "srio_pl_asymmetry_rcv_x2mr_x2rec_x2rn_x2rec_are_ari_test.sv"
`include "srio_pl_asymmetry_rcv_x1mr_x1rec_x1rn_x1rec_are_ari_test.sv"
`include "srio_pl_cw_retrain_timeout_lane2_test.sv"  
`include "srio_pl_cw_retrain_timeout_lanes4_test.sv" 
`include "srio_pl_cw_retrain_timeout_lanes8_test.sv"  
`include "srio_pl_cw_retrain_timeout_lanes16_test.sv" 
`include "srio_pl_cw_retrain_trnd_ret0_ret_fail_test.sv" 
`include "srio_pl_cw_retrain_trnd_ret1_ret_fail_test.sv" 
`include "srio_pl_asymmetry_x2mx_sx1mx_sx1mx2_sx1mx3_xwn_x2mx_test.sv"
`include "srio_pl_asymmetry_x2mx_sx1mx_sx1mx1_sx1mx2_axe_axi_test.sv"
`include "srio_pl_asymmetry_x1mx_x1mxa_test.sv"
`include "srio_pl_asymmetry_x2mx_x2mxa_test.sv"
`include "srio_pl_cw_retrain_timeout_1_test.sv"
`include "srio_pl_cw_retrain_timeout_retrain5_lanes16_test.sv"
`include "srio_pl_cw_retrain_retrain5_lanes16_test.sv"
`include "srio_pl_cw_retrain_retrain4_timeout_lanes8_test.sv" 
`include "srio_pl_cw_retrain_retrain5_lanes8_test.sv"
`include "srio_pl_cw_retrain_retrain5_timeout_lanes8_test.sv"
`include "srio_pl_cw_retrain_trnd_ret2_ret_fail_test.sv"  
`include "srio_pl_cw_retrain_retrain5_lanes2_test.sv"
`include "srio_pl_cw_retrain_retrain5_lanes4_test.sv"
`include "srio_pl_cw_retrain_retrain5_timeout_lanes4_test.sv"
`include "srio_pl_asymmetry_1x_port_req_test.sv"
`include "srio_pl_asymmetry_2x_port_req_test.sv"
`include "srio_pl_asymmetry_4x_port_req_test.sv"
`include "srio_pl_asymmetry_8x_port_req_test.sv"
`include "srio_pl_asymmetry_16x_port_req_test.sv"
`include "srio_pl_pkt_retry_cs_reset_test.sv"
`include "srio_pl_pkt_retry_cs_ors_reset_test.sv"
`include "srio_ll_lfc_vc_random_test.sv"
`include "srio_pl_cw_retrain_keep_alive_ret0_lanes2_test.sv"
`include "srio_pl_cw_retrain_keep_alive_ret0_lanes4_test.sv"
`include "srio_pl_cw_retrain_keep_alive_ret0_lanes8_test.sv"
`include "srio_pl_cw_retrain_keep_alive_ret0_lanes16_test.sv"
`include "srio_pl_cw_retrain_keep_alive_ret0_lanes1_test.sv"
`include "srio_ll_vc8_nwrite_swrite_test.sv"
`include "srio_ll_vc4_nwrite_swrite_test.sv"
`include "srio_ll_vc2_nwrite_swrite_test.sv"
`include "srio_pl_random_acc_gen_kind_test.sv"
`include "srio_pl_ies_oes_force_reinit_err_test.sv"
`include "srio_pl_force_1xmode_lane0_nx_support_test.sv"
`include "srio_pl_force_1xmode_lane0_2x_nx_support_test.sv"
`include "srio_pl_force_1xmode_laner_2x_support_test.sv"
`include "srio_pl_force_1xmode_laner_nx_support_test.sv"
`include "srio_pl_force_1xmode_laner_2x_nx_support_test.sv"
`include "srio_pl_cw_retrain_retrain5_timeout_lane1_test.sv"
`include "srio_pl_lane4_force_1x_mode_pa_na_test.sv"
`include "srio_pl_lane4_force_1x_mode_pa_retry_test.sv"
`include "srio_pl_lane4_force_1x_mode_laneR_pa_na_test.sv"
`include "srio_pl_lane4_force_1x_mode_laneR_pa_retry_test.sv"
`include "srio_pl_lane2_force_1x_mode_laneR_pa_na_test.sv"
`include "srio_pl_lane2_force_1x_mode_laneR_pa_retry_test.sv"
`include "srio_pl_timestamp_seq_err_test.sv"
`include "srio_ll_default_reset_test.sv"
`include "srio_ll_default_pa_na_reset_test.sv"
`include "srio_ll_default_pa_retry_reset_test.sv"
`include "srio_pl_delayed_pkt_acc_cs_test.sv"
`include "srio_pl_delayed_pkt_acc_retry_cs_test.sv"
`include "srio_pl_pa_cs_seq_ackid_test.sv"
`include "srio_pl_retry_pnack_cs_test.sv"
`include "srio_ll_nread_req_rand_resp_payload_test.sv"
`include "srio_ll_default_pa_na_b2b_test.sv"
`include "srio_ll_default_pa_retry_b2b_test.sv"
`include "srio_ll_default_pa_na_retry_b2b_test.sv"
`include "srio_ll_default_random_acc_pa_na_b2b_test.sv"
`include "srio_ll_default_random_acc_pa_retry_b2b_test.sv"
`include "srio_ll_default_random_acc_pa_b2b_test.sv"
`include "srio_ll_default_random_acc_pa_na_retry_b2b_test.sv"
`include "srio_pl_rfr_crc_corrupt_test.sv"
`include "srio_pl_rfr_to_pnack_corrupt_test.sv"
`include "srio_ll_resp_pkt_dis_test.sv"
`include "srio_ll_resp_payload_print_test.sv"
`include "srio_ll_resp_pri_error_test.sv"
`include "srio_pl_pkt_na_ackid_err_cs_test.sv"
`include "srio_pl_pkt_na_crc_err_cs_test.sv"
`include "srio_pl_pkt_na_non_maintenace_rep_stop_cs_test.sv"
`include "srio_pl_pkt_na_invalid_char_cs_test.sv"
`include "srio_pl_pkt_na_lack_buf_res_cs_test.sv"
`include "srio_pl_pkt_na_loss_descr_sync_cs_test.sv"
`include "srio_ll_ds_env1_env2_test.sv"
`include "srio_pl_pkt_prob_test.sv"
`include "srio_ll_nwrite_max_pkt_size_256b_test.sv"
`include "srio_ll_nread_req_link_init_test.sv"
`include "srio_ll_seq_order_pri_crf_retry_test.sv"
`endif
`include "srio_pl_pkt_early_final_crc_error_test.sv"
`include "srio_pl_gen3_incorrect_skip_ordered_lane_check_corrupt_test.sv"
`include "srio_pl_gen3_incorrect_skip_order_1_seq_test.sv"
`include "srio_pl_gen3_incorrect_skip_order_2_seq_test.sv"
`include "srio_pl_gen3_incorrect_skip_order_seq_test.sv"
`include "srio_pl_idle2_cs_marker_corrupt_test.sv"
`include "srio_pl_dis_nxmode_test.sv"
`include "srio_pl_nxmode_dis_test.sv"
`include "srio_pl_2xmode_1xmode_ln0_test.sv"
`include "srio_pl_2xmode_1xmode_ln1_test.sv"
`include "srio_ll_maintenance_rd_req_base_test.sv"
`include "srio_ll_msg_mseg_req_test.sv"
`include "srio_ll_msg_sseg_req_test.sv"
`include "srio_ll_gsm_dkill_home_test.sv"
`include "srio_ll_gsm_castout_test.sv"
`include "srio_ll_gsm_dkill_sharer_test.sv"
`include "srio_ll_gsm_flush_with_data_test.sv"
`include "srio_ll_gsm_flush_without_data_test.sv"
`include "srio_ll_gsm_ikill_home_test.sv"
`include "srio_ll_gsm_ikill_sharer_test.sv"
`include "srio_ll_gsm_io_read_home_test.sv"
`include "srio_ll_gsm_io_rd_owner_test.sv"
`include "srio_ll_gsm_iread_home_test.sv"
`include "srio_ll_gsm_rd_home_test.sv"
`include "srio_ll_gsm_rd_owner_test.sv"
`include "srio_ll_gsm_rd_to_own_home_test.sv"
`include "srio_ll_gsm_rd_to_own_owner_test.sv"
`include "srio_ll_gsm_tlbie_test.sv"
`include "srio_ll_gsm_tlbsync_test.sv"
`include "srio_ll_gsm_random_test.sv"
`include "srio_ll_callback_test.sv"
`include "srio_tl_callback_test.sv"
`include "srio_pl_callback_test.sv"
`include "srio_ll_ftype_error_test.sv"
`include "srio_ll_ttype_error_test.sv"
`include "srio_ll_max_size_error_test.sv"
`include "srio_ll_payload_error_test.sv"
`include "srio_ll_size_error_test.sv"
`include "srio_ll_no_payload_error_test.sv"
`include "srio_ll_no_payload_error_demote_test.sv"
`include "srio_ll_payload_exist_error_test.sv"
`include "srio_ll_atomic_compare_and_swap_error_test.sv"
`include "srio_ll_atomic_swap_error_test.sv"
`include "srio_ll_atomic_test_and_swap_payload_error_test.sv"
`include "srio_ll_doubleword_align_error_test.sv"
`include "srio_ll_msg_ssize_error_test.sv"
`include "srio_ll_msgseg_error_test.sv"
`include "srio_tl_destid_corrupt_callback_test.sv"
`include "srio_ll_resp_rsvd_sts_error_test.sv"
`include "srio_ll_resp_payload_error_test.sv"
`include "srio_pl_pkt_early_crc_error_test.sv"
`include "srio_pl_pkt_final_crc_error_test.sv"
`include "srio_pl_pkt_ackid_error_test.sv" 
`include "srio_pl_pkt_illegal_prio_error_test.sv" 
`include "srio_pl_pkt_illegal_crf_error_test.sv" 
`include "srio_pl_idle2_csfield_corruption_test.sv"
`include "srio_pl_idle2_psr_corruption_test.sv"
`include "srio_pl_idle2_csmarker_corruption_test.sv"
`include "srio_pl_idle2_desc_sync_break_corruption_test.sv"
`include "srio_ll_msg_interleaved_req_test.sv"
`include "srio_ll_io_random_test.sv"
`include "srio_ll_random_interleaved_test.sv"
`include "srio_ll_random_interleaved_weight_round_robin_test.sv"
`include "srio_ll_all_atomic_req_test.sv"
`include "srio_pl_nx_mode_support_disable_test.sv"
`include "srio_pl_2x_mode_support_disable_test.sv"
`include "srio_ll_read_write_test.sv"
`include "srio_ll_io_concurrent_trans.sv"
`include "srio_ll_msg_concurrent_req_test.sv"
`include "srio_ll_maintenance_wr_rd_test.sv"
`include "srio_ll_io_message_req_test.sv"
`include "srio_ll_io_message_doorbell_req_test.sv"
`include "srio_ll_unsupported_scr_dest_err_test.sv"
`include "srio_ll_nwrite_nread_34_addr_test.sv"
`include "srio_ll_nwrite_nread_50_addr_test.sv"
`include "srio_ll_nwrite_nread_66_addr_test.sv"
`include "srio_ll_parallel_mode_test.sv"
`include "srio_tl_pkt_tt_test.sv"
`include "srio_pl_nwrite_swrite_req_test.sv"
`include "srio_ll_illegal_io_trans_dec_test.sv"
`include "srio_ll_illegal_msg_trans_dec_test.sv"
`include "srio_ll_illegal_gsm_trans_dec_test.sv"
`include "srio_ll_ds_concurrent_test.sv"
`include "srio_ll_ds_max_seg_support_test.sv"
`include "srio_ll_ds_mtu_reserved_test.sv"
`include "srio_ll_ds_s_e_err_test.sv"
`include "srio_ll_multi_vc_nwrite_swrite_test.sv"
`include "srio_ll_traffic_mgmt_tm_type_mode_err_test.sv"
`include "srio_ll_maintenance_ds_test.sv"
`include "srio_ll_ds_traffic_mgmt_diff_operation_test.sv"
`include "srio_ll_lfc_pri_error_test.sv"
`include "srio_ll_lfc_xoff_test.sv"
`include "srio_ll_lfc_xon_test.sv"
`include "srio_ll_msg_interleaved_out_of_order_test.sv"
`include "srio_ll_msg_mseg_req_with_msgseg_err_test.sv"
`include "srio_ll_msg_mseg_req_with_msglen_err_test.sv"
`include "srio_ll_msg_mseg_req_max_pld_test.sv"
`include "srio_ll_msg_mseg_req_with_sseg_neqt_ssize_err_test.sv"
`include "srio_ll_msg_mseg_req_with_cseg_neqt_ssize_err_test.sv"
`include "srio_ll_msg_mseg_req_with_eseg_gt_ssize_err_test.sv"
`include "srio_ll_msg_mseg_req_without_payload_err_test.sv"
`include "srio_ll_atomic_invalid_size.sv"
`include "srio_ll_msg_mseg_req_with_lastseg_err_test.sv"
`include "srio_tl_invalid_tt_callback_test.sv"
`include "srio_ll_msg_unsupported_trans_test.sv"
`include "srio_ll_db_unsupported_trans_test.sv"
`include "srio_ll_illegal_ftpe_ttype_callback_test.sv"
`include "srio_ll_msg_max_pld_with_mbox_letter_test.sv"
`include "srio_pl_nxmode_sl_test.sv"
`include "srio_ll_msg_cov_test.sv"
`include "srio_ll_io_gsm_less_payload_test.sv"
`include "srio_pl_crc32_err_cb_test.sv"
`include "srio_pl_cg_invalid_for_skip_cb_test.sv"
`include "srio_pl_sop_padded_length_not8multiple_test.sv"
`include "srio_pl_gen3_incorrect_spacing_cw_bw_sc_cw_test.sv"
`include "srio_pl_sync_reset_s_to_ns_test.sv"
`include "srio_pl_aet_test.sv"
`include "srio_pl_aet_tplus_hold_test.sv"
`include "srio_pl_aet_tplus_tincr_test.sv"
`include "srio_pl_aet_tplus_tdecr_test.sv"
`include "srio_pl_aet_tminus_hold_incr_test.sv"
`include "srio_pl_aet_tminus_incr_incr_test.sv"
`include "srio_pl_aet_tminus_incr_decr_test.sv"
`include "srio_pl_aet_tminus_incr_hold_test.sv"
`include "srio_pl_aet_tminus_hold_decr_test.sv"
`include "srio_pl_aet_tminus_test.sv"
`include "srio_pl_aet_tplus_random_test.sv"
`include "srio_pl_aet_tminus_random_test.sv"
`include "srio_pl_aet_preset_test.sv"
`include "srio_pl_aet_rst_test.sv"
`include "srio_pl_aet_not_supported_err_test.sv"
`include "srio_pl_idle2_cs_field_aet_cmd_corrupt_cb_test.sv"
`include "srio_pl_idle2_cs_field_aet_ack_nack_corrupt_cb_test.sv"
`include "srio_pl_idle2_mmmm_seq_corruption_test.sv"
`include "srio_pl_idle2_KR_seq_corruption_test.sv"
`include "srio_pl_idle2_cg_between_clk_comp_check_err_test.sv"
`include "srio_pl_idle2_MDDDD_sync_sequence_corrupt_err_test.sv"
`include "srio_pl_idle2_invalid_MDDDD_sync_seq_err_test.sv" 
`include "srio_pl_dis_2xmode_test.sv"
`include "srio_pl_dis_1xmode_ln0_test.sv"
`include "srio_pl_dis_1xmode_ln1_test.sv"
`include "srio_pl_dis_1xmode_ln2_test.sv"
`include "srio_pl_dis_sl_test.sv"
`include "srio_pl_2xmode_sl_test.sv"
`include "srio_pl_sync_reset_ns3_to_ns_test.sv"
`include "srio_pl_sync_reset_ns1_to_ns_test.sv"
`include "srio_pl_2xmode_2x_rec_test.sv"
`include "srio_pl_1xmode_ln0_sl_test.sv"
`include "srio_pl_1xmode_ln0_1x_rec_test.sv"
`include "srio_pl_1xmode_ln1_sl_test.sv"
`include "srio_pl_1xmode_ln1_1x_rec_test.sv"
`include "srio_pl_1xmode_ln2_sl_test.sv"
`include "srio_pl_1xmode_ln2_1x_rec_test.sv"
`include "srio_pl_2x_rec_2xmode_test.sv"
`include "srio_pl_2x_rec_1xmode_ln0_test.sv"
`include "srio_pl_2x_rec_1xmode_ln1_test.sv"
`include "srio_pl_2x_rec_sl_test.sv"
`include "srio_pl_1x_rec_sl_test.sv"
`include "srio_pl_1x_rec_1xmode_ln0_test.sv"
`include "srio_pl_1x_rec_1xmode_ln1_test.sv"
`include "srio_pl_1x_rec_1xmode_ln2_test.sv"
`include "srio_pl_nxm_dis_sl_test.sv"  
`include "srio_pl_nxm_dis_1xm0_test.sv" 
`include "srio_pl_nxm_dis_1xm1_test.sv" 
`include "srio_pl_nxm_dis_1xm2_test.sv" 
`include "srio_pl_nxm_dis_2xm_test.sv"
`include "srio_pl_nxm_dis_nxm_test.sv"
`include "srio_pl_x1m1_x1r_sl_test.sv"
`include "srio_pl_x1m2_x1r_sl_test.sv"
`include "srio_pl_reset_seek_test.sv"
`include "srio_pl_reset_discovery_test.sv"
`include "srio_pl_reset_nx_mode_test.sv"
`include "srio_pl_reset_2xmode_test.sv"
`include "srio_pl_reset_nx_recovery_test.sv"
`include "srio_pl_reset_2x_recovery_test.sv"
`include "srio_pl_reset_1xmode_ln0_test.sv"
`include "srio_pl_reset_1xmode_ln1_test.sv"
`include "srio_pl_reset_1xmode_ln2_test.sv"
`include "srio_pl_reset_1xmode_recovery_test.sv"
`include "srio_pl_force_reinit_discovery_test.sv" 
`include "srio_pl_force_reinit_seek_test.sv"
`include "srio_pl_force_reinit_2xmode_test.sv"
`include "srio_pl_force_reinit_nx_mode_test.sv"
`include "srio_pl_force_reinit_2x_recovery_test.sv"
`include "srio_pl_force_reinit_1xmode_ln0_test.sv"
`include "srio_pl_force_reinit_1xmode_ln1_test.sv"
`include "srio_pl_force_reinit_1xmode_ln2_test.sv"
`include "srio_pl_force_reinit_1xmode_recovery_test.sv"
`include "srio_pl_force_reinit_test.sv"
`include "srio_pl_link_req_rst_3_b2b_sop_link_req_rst_cs_test.sv"
`include "srio_pl_link_req_rst_2_b2b_sop_2_b2b_link_req_rst_cs_test.sv"
`include "srio_pl_trans_scramble_enable_test.sv"
`include "srio_pl_diff_idle_sel_test.sv"
`include "srio_pl_skew_max_min_test.sv"
`include "srio_pl_gen2_a1_a2_a2_sm_test.sv"
`include "srio_pl_align_error_test.sv"
`include "srio_ll_invalid_tt_test.sv"
`include "srio_pl_nop_cs_test.sv"
`include "srio_pl_sop_cs_test.sv"
`include "srio_pl_eop_cs_test.sv"
`include "srio_pl_link_req_input_dev_cs_test.sv"
`include "srio_pl_link_req_rst_dev_cs_test.sv"
`include "srio_pl_restart_rty_cs_test.sv"
`include "srio_pl_stomp_cs_test.sv"
`include "srio_pl_align_reset_sm_test.sv" 
`include "srio_pl_sop_nwrite_eop_test.sv"
`include "srio_pl_sync_break_all_lanes_test.sv"
`include "srio_pl_ns1_ns2_ns1_ns2_sm_all_lanes_test.sv"
`include "srio_pl_ns1_ns2_ns_sm_all_lanes_test.sv"
`include "srio_pl_sync_sm_all_lanes_test.sv"
`include "srio_pl_ns1_ns2_ns3_ns2_ns_sm_all_lanes_test.sv"
`include "srio_pl_ns1_ns2_ns3_ns2_ns1_sm_all_lanes_test.sv"
`include "srio_pl_link_req_rst_4_b2b_cs_test.sv"
`include "srio_pl_link_req_rst_3_b2b_status_cs_link_req_rst_test.sv"
`include "srio_pl_link_req_rst_3_b2b_non_status_cs_link_req_rst_test.sv"
`include "srio_pl_link_req_rst_2_b2b_non_status_cs_2_link_req_rst_test.sv"
`include "srio_pl_link_req_rst_1_b2b_non_status_cs_3_link_req_rst_test.sv"
`include "srio_pl_link_req_rst_1_b2b_status_cs_3_link_req_rst_test.sv"
`include "srio_pl_link_req_rst_2_b2b_status_cs_2_link_req_rst_test.sv"
`include "srio_pl_link_req_rst_b2b_status_cs_link_req_rst_test.sv"
`include "srio_pl_link_req_rst_port_4_b2b_cs_test.sv"
`include "srio_pl_link_req_rst_port_3_b2b_status_cs_link_req_rst_port_test.sv"
`include "srio_pl_link_req_rst_port_3_b2b_non_status_cs_link_req_rst_port_test.sv"
`include "srio_pl_link_req_rst_port_2_b2b_non_status_cs_2_link_req_rst_port_test.sv"
`include "srio_pl_link_req_rst_port_1_b2b_status_cs_3_link_req_rst_port_test.sv"
`include "srio_pl_link_req_rst_port_1_b2b_non_status_cs_3_link_req_rst_port_test.sv"
`include "srio_pl_link_req_rst_port_2_b2b_status_cs_2_link_req_rst_port_test.sv"
`include "srio_pl_link_req_rst_port_b2b_status_cs_link_req_rst_port_test.sv"
`include "srio_pl_reset_a1_na_a_test.sv"
`include "srio_pl_reset_a2_na_a_test.sv"
`include "srio_pl_reset_a3_na_a_test.sv"
`include "srio_pl_sync_signal_detect_ns1_ns_test.sv"
`include "srio_pl_sync_signal_detect_ns3_ns_test.sv"
`include "srio_pl_sync_signal_detect_s_ns_test.sv"
`include "srio_pl_sync_signal_detect_s1_ns_test.sv"
`include "srio_pl_sync_signal_detect_s3_ns_test.sv"
`include "srio_pl_sync_signal_detect_s4_ns_test.sv"
`include "srio_pl_sync_reset_s1_to_ns_test.sv" 
`include "srio_pl_sync_reset_s3_to_ns_test.sv" 
`include "srio_pl_sync_reset_s4_to_ns_test.sv"
`include "srio_pl_nxm_nxr_nxrn_nxm_test.sv" //GEN3
`include "srio_pl_nxm_nxr_nxrn_2x_test.sv"
`include "srio_pl_nxm_nxr_nxrn_x1m0_test.sv"
`include "srio_pl_nxm_nxr_nxrn_x1m1_test.sv"
`include "srio_pl_nxm_nxr_nxrn_x1m2_test.sv"
`include "srio_pl_x2m_x2r_x2rn_x2r_x2m_test.sv"
`include "srio_pl_x2m_x2r_x2rn_x2r_x1m0_test.sv"
`include "srio_pl_x2m_x2r_x2rn_x2r_x1m1_test.sv"
`include "srio_pl_x1m0_x1r_x1rn_x1r_x1m0_test.sv"
`include "srio_pl_x1m1_x1r_x1rn_x1r_x1m1_test.sv"
`include "srio_pl_x1m2_x1r_x1rn_x1r_x1m2_test.sv"
`include "srio_pl_nxr_nxrn_nxr_sil_test.sv"
`include "srio_pl_x1m0_x1r_x1rn_x1r_sl_test.sv"
`include "srio_pl_x1m1_x1r_x1rn_x1r_sl_test.sv"
`include "srio_pl_x1m2_x1r_x1rn_x1r_sl_test.sv"
`include "srio_pl_x2m_x2r_x2rn_x2r_sil_test.sv"
`include "srio_pl_force_reinit_nxretrain_test.sv"
`include "srio_pl_force_reinit_2xretrain_test.sv"
`include "srio_pl_force_reinit_1xretrain_test.sv"
`include "srio_pl_reset_nxretrain_test.sv"
`include "srio_pl_reset_2xretrain_test.sv"
`include "srio_pl_reset_1xretrain_test.sv"
`include "srio_pl_nxm_nxr_test.sv"
`include "srio_pl_nxr_nxm_test.sv" 
`include "srio_pl_nxr_1xm0_test.sv"  
`include "srio_pl_nxr_1xm1_test.sv"
`include "srio_pl_nxr_1xm2_test.sv"
`include "srio_pl_nxr_sil_test.sv"
`include "srio_pl_nxr_2xm_test.sv"
`include "srio_pl_force_reinit_nx_recovery_test.sv"
`include "srio_pl_sop_with_eop_cs_test.sv"
`include "srio_pl_sop_stomp_cs_test.sv"
`include "srio_pl_sop_link_req_cs_test.sv"
`include "srio_pl_sop_link_req_rst_cs_test.sv"
`include "srio_pl_link_response_cs_test.sv"
`include "srio_pl_gen3_a_a2_a3_a4_sm_test.sv"
`include "srio_pl_gen3_a3_a4_a5_a3_sm_test.sv" 
`include "srio_pl_gen3_a3_a4_a6_a3_sm_test.sv"  
`include "srio_pl_gen3_ns2_ns3_ns1_sm_all_lanes_test.sv"
`include "srio_pl_sop_link_req_inp_stat_callback_test.sv"
`include "srio_pl_sop_restart_rty_callback_test.sv"
`include "srio_pl_sop_link_req_rst_dev_callback_test.sv"
`include "srio_pl_gen3_sop_eop_padded_cs_test.sv"
`include "srio_pl_gen3_eop_padded_cs_test.sv"
`include "srio_pl_gen3_reset_na2_na_test.sv"
`include "srio_pl_gen3_reset_na3_na_test.sv"
`include "srio_pl_gen3_reset_na1_na_test.sv"
`include "srio_pl_gen3_reset_a_na_test.sv"
`include "srio_pl_gen3_reset_a3_na_test.sv"
`include "srio_pl_gen3_reset_a4_na_test.sv"
`include "srio_pl_gen3_reset_a5_na_test.sv"
`include "srio_pl_gen3_reset_a7_na_test.sv"
`include "srio_pl_gen3_reset_a6_na_test.sv"
`include "srio_pl_gen3_reset_a1_na_test.sv"
`include "srio_pl_gen3_reset_a2_na_test.sv"
`include "srio_pl_gen3_reset_ns3_ns_test.sv"
`include "srio_pl_gen3_reset_ns4_ns_test.sv"
`include "srio_pl_gen3_reset_s_ns_test.sv"
`include "srio_pl_gen3_reset_s1_ns_test.sv"
`include "srio_pl_gen3_reset_s2_ns_test.sv"
`include "srio_pl_gen3_reset_ns1_ns_test.sv"
`include "srio_pl_start_cw_open_context_err_test.sv"
`include "srio_pl_end_cw_closed_context_err_test.sv"
`include "srio_pl_end_cw_corrupted_to_data_err_test.sv"
`include "srio_pl_gen3_incorrect_skip_marker_fixed_value_cb_test.sv"
`include "srio_pl_gen3_incorrect_lc_flwd_by_sc_cw_test.sv"
`include "srio_pl_aligned_aligned1_notaligned_sm_test.sv"
`include "srio_pl_lane_align_sm_test.sv"
`include "srio_pl_cs_insertion_cb_test.sv"
`include "srio_pl_lane_data_cntl_corruption_test.sv"
`include "srio_pl_idle2_krrr_insert_sequence_cb_test.sv"
`include "srio_pl_pkt_crc_corruption_test.sv"
`include "srio_pl_cs_crc_corrupt_test.sv"
`include "srio_gen3_pkt_crc_cb_corrupt_test.sv"
`include "srio_pl_sop_idle2_eop_test.sv"
`include "srio_pl_sop_idle2_lreq_test.sv"
`include "srio_ll_port_resp_timeout_reg_test.sv" 
`include "srio_tl_ds_scrid_err_cb_test.sv"
`include "srio_ll_db_pkt_ratio_test.sv"
`include "srio_ll_io_pkt_ratio_test.sv"
`include "srio_ll_gsm_pkt_ratio_test.sv"
`include "srio_ll_msg_pkt_ratio_test.sv"
`include "srio_ll_nwrite_nread_mem_access_test.sv"
`include "srio_ll_ds_corner_case_total_pkt_80byte_test.sv" 
`include "srio_ll_ds_interleaved_test.sv"
`include "srio_ll_ds_mseg_single_mtu_test.sv"
`include "srio_ll_ds_pkt_ratio_test.sv"
`include "srio_ll_ds_traffic_mgmt_random_basic_stream_test.sv"
`include "srio_ll_ds_traffic_mgmt_random_rate_stream_test.sv"
`include "srio_ll_ds_traffic_mgmt_random_credit_stream_test.sv"
`include "srio_ll_vc_ds_mseg_req_test.sv"
`include "srio_ll_ds_mseg_req_with_sseg_neqt_mtu_err_test.sv"
`include "srio_ll_ds_mseg_req_with_cseg_neqt_mtu_err_test.sv"
`include "srio_ll_ds_mseg_req_without_payload_err_test.sv"
`include "srio_ll_ds_mseg_req_with_invalid_pdulen_err_test.sv"
`include "srio_ll_ds_max_pdu_streamid_test.sv"
`include "srio_ll_traffic_mgmt_random_test.sv"
`include "srio_ll_ds_mtu_error_test.sv" 
`include "srio_ll_ds_pdu_error_test.sv"
`include "srio_ll_ds_sop_error_test.sv"
`include "srio_ll_ds_eop_error_test.sv"
`include "srio_ll_ds_pad_error_test.sv"
`include "srio_ll_ds_odd_error_test.sv"
`include "srio_ll_ds_sseg_req_test.sv"
`include "srio_ll_ds_mseg_req_test.sv"
`include "srio_ll_ds_max_min_pdu_mtu_test.sv"
`include "srio_ll_ds_traffic_mgmt_basic_stream_test.sv"
`include "srio_ll_ds_traffic_mgmt_rate_control_test.sv"
`include "srio_ll_ds_traffic_mgmt_credit_control_test.sv"
`include "srio_ll_ds_traffic_mgmt_credit_rate_control_test.sv"
`include "srio_ll_ds_pdu_length_err_test.sv"
`include "srio_ll_ds_normal_error_test.sv"
`include "srio_ll_io_ds_test.sv"
`include "srio_ll_ds_traffic_mgmt_mask_err_test.sv"
`include "srio_ll_atomic_req_followedby_any_req_err_test.sv"
`include "srio_ll_io_random_with_speci_src_tid_test.sv"
`include "srio_ll_io_random_with_speci_src_tid_same_sc_des_err_test.sv"
`include "srio_ll_msg_with_same_mbox_letter_test.sv"
`include "srio_ll_msg_with_same_mbox_letter_scid_desid_err_test.sv"
`include "srio_ll_ds_mseg_with_speci_cos_req_test.sv"
`include "srio_ll_ds_mseg_with_speci_cos_scid_desid_err_req_test.sv"
`include "srio_pl_pkt_acc_cs_test.sv"
`include "srio_pl_seek_1xmode_ln0_test.sv" 
`include "srio_pl_seek_1xmode_ln2_test.sv" 
`include "srio_pl_sync_break_test.sv"
`include "srio_pl_sync_sm_test.sv"
`include "srio_pl_clck_comp_code_group_cs_test.sv"
`include "srio_pl_asymmetry_silent_test.sv"
`include "srio_pl_nxm_asymetry_test.sv"
`include "srio_pl_2xm_asymmetry_test.sv"  
`include "srio_pl_reset_asymmetry_test.sv" 
`include "srio_pl_force_reinit_asymmetry_test.sv"
`include "srio_pl_ns1_ns2_ns3_ns2_ns_sm_test.sv"
`include "srio_pl_ns1_ns2_ns3_ns2_ns1_sm_test.sv"
`include "srio_pl_gen3_ns2_ns3_ns1_sm_test.sv"
`include "srio_pl_env1_sop_link_req_env2_disabled_test.sv" 
`include "srio_pl_env1_sop_link_req_rst_dev_env2_disabled_test.sv"
`include "srio_pl_env1_sop_stomp_env2_disabled_test.sv" 
`include "srio_pl_env1_sop_restart_rty_env2_disabled_test.sv"
`include "srio_pl_env1_sop_eop_env2_disabled_test.sv" 
`include "srio_pl_sop_stomp_callback_test.sv" 
`include "srio_pl_reset_na2_na_test.sv"
`include "srio_pl_reset_na1_na_test.sv"
`include "srio_pl_align_error_2_sm_test.sv"
`include "srio_pl_retrain_disable_test.sv"
`include "srio_pl_idle2_seq_with_status_control_cs_err_test.sv"
`include "srio_pl_corrupt_eop_stomp_test.sv"
`include "srio_ll_multiple_ack_default_test.sv"
`include "srio_ll_multiple_ack_with_pa_retry_ratio_default_test.sv"
`include "srio_ll_multiple_ack_with_pa_na_ratio_default_test.sv"
`include "srio_ll_default_pa_na_test.sv"
`include "srio_ll_default_pa_retry_test.sv"
`include "srio_ll_default_random_acc_pa_na_test.sv"
`include "srio_ll_default_random_acc_pa_retry_test.sv"
`include "srio_ll_default_random_acc_pa_test.sv"
`include "srio_ll_default_max_random_acc_pa_retry_test.sv"
`include "srio_ll_default_max_random_acc_pa_test.sv"
`include "srio_ll_default_max_random_acc_pa_na_test.sv" 
`include "srio_ll_default_pa_na_retry_test.sv"
`include "srio_pl_cw_train_incr_tap0_test.sv"
`include "srio_pl_cw_train_decr_tap0_test.sv"
`include "srio_pl_cw_train_incr_decr_tap0_test.sv"
`include "srio_pl_cw_train_kind_disabled_test.sv"
`include "srio_pl_cw_train_hold_test.sv"
`include "srio_pl_cw_train_initialize_test.sv"
`include "srio_pl_cw_train_preset_random_test.sv"
`include "srio_pl_cw_train_initialize_random_test.sv"
`include "srio_pl_cw_train_hold_random_test.sv"
`include "srio_pl_cw_train_incr_random_test.sv"
`include "srio_pl_cw_train_decr_random_test.sv"
`include "srio_pl_cw_train1_cw_train_fail_test.sv"
`include "srio_pl_dme_test.sv"
`include "srio_pl_dme_hold_test.sv"
`include "srio_pl_dme_decr_test.sv"
`include "srio_pl_dme_incre_test.sv"
`include "srio_pl_dme_init_test.sv"
`include "srio_pl_dme_prst_test.sv"
`include "srio_pl_dme_max_limit_test.sv"
`include "srio_pl_dme1_dmef_test.sv"
`include "srio_pl_dme1_to_untrk_dmet2_test.sv"
`include "srio_pl_ackid_status_corrupt_err_test.sv"
`include "srio_pl_pnack_diff_cause_gen1_err_test.sv"
`include "srio_pl_pnack_diff_cause_gen2_err_test.sv"
`include "srio_pl_pnack_diff_cause_gen3_err_test.sv"
`include "srio_ll_nwrite_max_byte_err_test.sv"
`include "srio_pl_gen3_cwl_descr_seed_skip_order_corrupt_test.sv"
`include "srio_pl_gen3_sync_break_test.sv"
`include "srio_pl_gen3_sync_sm_s_s1_s2_all_lanes_test.sv"
`include "srio_pl_gen3_sync_sm_s_s1_s2_test.sv"
`include "srio_pl_only_idle_no_pkt_test.sv"
`include "srio_ll_nwrite_80bytes_less_greater_test.sv"
`include "srio_pl_gen3_cwl_descr_seed_skip_order_rand_corrupt_test.sv"
endpackage :srio_test_lib_pkg
