////////////////////////////////////////////////////////////////////////////////
//(c) Copyright 2013 Mobiveil, Inc. All rights reserved
//
// File    :  srio_pl_callback.sv
// Project :  srio vip
// Purpose :  Physical Layer Call Back
// Author  :  Mobiveil
//
// Physical Layer Callback class.
//
//////////////////////////////////////////////////////////////////////////////// 
typedef class srio_pl_data_trans;

class srio_pl_callback extends uvm_callback; 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : New
/// Description : Constructor method for srio_pl_callback class.
///////////////////////////////////////////////////////////////////////////////////////////////
function new (string name = "srio_pl_callback"); 
super.new(name); 

endfunction 

static string type_name = "srio_pl_callback"; 		///< Class name declared as string. Returned when get_type_name is called.


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : get_type_name
/// Description : This method will return the class name when called.
///////////////////////////////////////////////////////////////////////////////////////////////
virtual function string get_type_name(); 
return type_name; 
endfunction



///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_trans_generated
/// Description : Callback method for trans generated on tx path.
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_trans_generated(ref srio_trans tx_srio_trans);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_trans_received
/// Description : Callback method for trans received on tx path.
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_trans_received(ref srio_trans rx_srio_trans);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane0
/// Description : Callback method for codegroup/codeword generated on lane driver instance '0'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane0(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config );
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane1
/// Description : Callback method for codegroup/codeword generated on lane driver instance '1'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane1(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane2
/// Description : Callback method for codegroup/codeword generated on lane driver instance '2'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane2(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane3
/// Description : Callback method for codegroup/codeword generated on lane driver instance '3'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane3(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane4
/// Description : Callback method for codegroup/codeword generated on lane driver instance '4'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane4(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane5
/// Description : Callback method for codegroup/codeword generated on lane driver instance '5'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane5(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane6
/// Description : Callback method for codegroup/codeword generated on lane driver instance '6'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane6(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane7
/// Description : Callback method for codegroup/codeword generated on lane driver instance '7'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane7(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane8
/// Description : Callback method for codegroup/codeword generated on lane driver instance '8'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane8(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane9
/// Description : Callback method for codegroup/codeword generated on lane driver instance '9'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane9(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane10
/// Description : Callback method for codegroup/codeword generated on lane driver instance '10'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane10(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane11
/// Description : Callback method for codegroup/codeword generated on lane driver instance '11'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane11(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane12
/// Description : Callback method for codegroup/codeword generated on lane driver instance '12'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane12(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane13
/// Description : Callback method for codegroup/codeword generated on lane driver instance '13'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane13(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane14
/// Description : Callback method for codegroup/codeword generated on lane driver instance '14'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane14(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_generated_lane15
/// Description : Callback method for codegroup/codeword generated on lane driver instance '15'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_generated_lane15(ref srio_pl_lane_data tx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane0
/// Description : Callback method for codegroup/codeword received on lane handler instance '0'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane0(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane1
/// Description : Callback method for codegroup/codeword received on lane handler instance '1'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane1(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane2
/// Description : Callback method for codegroup/codeword received on lane handler instance '2'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane2(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane3
/// Description : Callback method for codegroup/codeword received on lane handler instance '3'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane3(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane4
/// Description : Callback method for codegroup/codeword received on lane handler instance '4'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane4(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane5
/// Description : Callback method for codegroup/codeword received on lane handler instance '5'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane5(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane6
/// Description : Callback method for codegroup/codeword received on lane handler instance '6'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane6(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane7
/// Description : Callback method for codegroup/codeword received on lane handler instance '7'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane7(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane8
/// Description : Callback method for codegroup/codeword received on lane handler instance '8'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane8(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane9
/// Description : Callback method for codegroup/codeword received on lane handler instance '9'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane9(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane10
/// Description : Callback method for codegroup/codeword received on lane handler instance '10'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane10(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane11
/// Description : Callback method for codegroup/codeword received on lane handler instance '11'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane11(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane12
/// Description : Callback method for codegroup/codeword received on lane handler instance '12'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane12(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane13
/// Description : Callback method for codegroup/codeword received on lane handler instance '13'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane13(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane14
/// Description : Callback method for codegroup/codeword received on lane handler instance '14'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane14(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_cg_received_lane15
/// Description : Callback method for codegroup/codeword received on lane handler instance '15'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_cg_received_lane15(ref srio_pl_lane_data rx_srio_cg,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane0
/// Description : Callback method for idle2 cs field received on lane handler instance '0'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane0(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane1
/// Description : Callback method for idle2 cs field received on lane handler instance '1'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane1(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane2
/// Description : Callback method for idle2 cs field received on lane handler instance '2'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane2(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane3
/// Description : Callback method for idle2 cs field received on lane handler instance '3'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane3(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane4
/// Description : Callback method for idle2 cs field received on lane handler instance '4'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane4(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane5
/// Description : Callback method for idle2 cs field received on lane handler instance '5'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane5(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane6
/// Description : Callback method for idle2 cs field received on lane handler instance '6'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane6(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane7
/// Description : Callback method for idle2 cs field received on lane handler instance '7'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane7(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane8
/// Description : Callback method for idle2 cs field received on lane handler instance '8'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane8(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane9
/// Description : Callback method for idle2 cs field received on lane handler instance '9'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane9(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane10
/// Description : Callback method for idle2 cs field received on lane handler instance '10'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane10(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane11
/// Description : Callback method for idle2 cs field received on lane handler instance '11'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane11(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane12
/// Description : Callback method for idle2 cs field received on lane handler instance '12'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane12(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane13
/// Description : Callback method for idle2 cs field received on lane handler instance '13'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane13(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane14
/// Description : Callback method for idle2 cs field received on lane handler instance '14'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane14(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_aet_cs_received_lane15
/// Description : Callback method for idle2 cs field received on lane handler instance '15'
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_aet_cs_received_lane15(ref srio_pl_rcvd_cs_field_data rx_cs_fld);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_trans_transmit
/// Description : Callback method for Control Symbola and Packet to be transmitted
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_trans_transmit(ref srio_pl_data_trans tx_gen,srio_trans srio_trans_in);
endtask 

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane0
/// Description : Callback method for character transmitted on lane0
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane0(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask 


///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane1
/// Description : Callback method for character transmitted on lane1
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane1(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane2
/// Description : Callback method for character transmitted on lane2
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane2(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane3
/// Description : Callback method for character transmitted on lane3
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane3(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane4
/// Description : Callback method for character transmitted on lane4
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane4(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane5
/// Description : Callback method for character transmitted on lane5
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane5(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane6
/// Description : Callback method for character transmitted on lane6
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane6(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane7
/// Description : Callback method for character transmitted on lane7
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane7(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane8
/// Description : Callback method for character transmitted on lane65
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane8(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane9
/// Description : Callback method for character transmitted on lane9
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane9(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane10
/// Description : Callback method for character transmitted on lane10
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane10(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane11
/// Description : Callback method for character transmitted on lane11
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane11(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane12
/// Description : Callback method for character transmitted on lane12
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane12(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane13
/// Description : Callback method for character transmitted on lane13
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane13(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane14
/// Description : Callback method for character transmitted on lane14
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane14(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask

///////////////////////////////////////////////////////////////////////////////////////////////
/// Name : srio_pl_char_transmitted_lane15
/// Description : Callback method for character transmitted on lane15
///////////////////////////////////////////////////////////////////////////////////////////////
virtual task srio_pl_char_transmitted_lane15(ref bit [0:65] idle_field_char,srio_env_config env_config);
endtask
endclass : srio_pl_callback 

