////////////////////////////////////////////////////////////////////////////////
//(c) Copyright 2013 Mobiveil, Inc. All rights reserved
//
// File    : srio_pl_gen3_reset_ns3_ns_test .sv
// Project :  srio vip
// Purpose :  LANE ALIGN STATE MACHINE
// Author  :  Mobiveil
//
// // 1.wait for  NO_SYNC_3  .
// 2. apply reset.after that deassarted reset.
// 3. After state changes wait for NO_SYNC_3.
// 4.After link initialized,send nread packets.
// Supported by only  Gen3 mode
////////////////////////////////////////////////////////////////////////////////

class srio_pl_gen3_reset_ns3_ns_test extends srio_base_test;

  `uvm_component_utils(srio_pl_gen3_reset_ns3_ns_test)
   rand int num;
   srio_ll_nread_req_seq nread_req_seq;
   
  function new(string name, uvm_component parent=null);
    super.new(name, parent);
     endfunction
  
     task run_phase( uvm_phase phase );
    super.run_phase(phase);
      
    nread_req_seq = srio_ll_nread_req_seq::type_id::create("nread_req_seq");

     phase.raise_objection( this );
     num = $urandom_range(32'd2,32'd0); 
      if(env_config1.num_of_lanes == 1) begin //{ 
      case(num)  //{
      32'd0 : wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[num].current_sync_state == NO_SYNC_3);
      32'd1 : wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[num].current_sync_state == NO_SYNC_3);
      32'd2 : wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[num].current_sync_state == NO_SYNC_3);
      endcase //}
      end //} 
      else if(env_config1.num_of_lanes == 2) begin //{
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[0].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[1].current_sync_state == NO_SYNC_3);  
      end //}
      else if(env_config1.num_of_lanes == 4) begin //{
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[0].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[1].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[2].current_sync_state == NO_SYNC_3);  
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[3].current_sync_state == NO_SYNC_3);
        
      end //}
      else if(env_config1.num_of_lanes == 8) begin //{
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[0].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[1].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[2].current_sync_state == NO_SYNC_3);  
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[3].current_sync_state == NO_SYNC_3);  
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[4].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[5].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[6].current_sync_state == NO_SYNC_3);  
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[7].current_sync_state == NO_SYNC_3);  
      end //}
      else  begin //{
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[0].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[1].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[2].current_sync_state == NO_SYNC_3);  
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[3].current_sync_state == NO_SYNC_3);  
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[4].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[5].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[6].current_sync_state == NO_SYNC_3);  
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[7].current_sync_state == NO_SYNC_3);   
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[8].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[9].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[10].current_sync_state == NO_SYNC_3);  
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[11].current_sync_state == NO_SYNC_3);  
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[12].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[13].current_sync_state == NO_SYNC_3);
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[14].current_sync_state == NO_SYNC_3);  
      wait(env1.pl_agent.pl_monitor.rx_monitor.lane_handle_ins[15].current_sync_state == NO_SYNC_3);  
      end //}


      env1.pl_agent.pl_driver.srio_if.srio_rst_n = 0;
      #1000ns;
      env1.pl_agent.pl_driver.srio_if.srio_rst_n = 1;
      nread_req_seq.start(env1.e_virtual_sequencer);
      #2000ns;     
      phase.drop_objection(this);
    
  endtask

  
endclass


